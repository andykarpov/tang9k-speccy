--
--Written by GowinSynthesis
--Product Version "GowinSynthesis V1.9.8.05"
--Fri May 12 17:32:10 2023

--Source file index table:
--file0 "\/opt/Gowin/IDE/ipcore/PSRAM_HS/data/PSRAM_TOP.v"
--file1 "\/opt/Gowin/IDE/ipcore/PSRAM_HS/data/psram_code.v"
`protect begin_protected
`protect version="2.1"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.1"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2021-10",key_method="rsa"
`protect key_block
G1wBuWOXxf1xs6eG6+/gC5frKt3bDXAvtVl9OLT4Ixe5GHT5kBLXJthlfTTZK7+f0QQ5WeIXiL8n
FS0lTmuoiYpgmHVRdKwyHCvPOxV8BOK+f/2+kiyPo694hOArNgQVzDW8hioZUsDSuD38IXBHSgKy
6+7aXdlMVj/WDaCNzs9dmVKyYY5z6MFk5lEeZkXzMeHq8LrWXYGaaInwlL61L/WJS3CyOrbr2gpc
CEvtRtrLxnZzlSX4S2Kxff5FNdFl33OT9kK8MSwY/W7bIPHDgZDcQtANVI4OdknGpyUgV4T1Lss4
HnT9SHMZATy4UYVh1UasKsXXw1GHe8PdxPQk/A==

`protect encoding=(enctype="base64", line_length=76, bytes=326048)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cbc"
`protect data_block
Ud2M7XAthOq7fbZc4XZKKXaDv2aiQuDp6d5GsCGyFAwgilINKNNk2uHoqhdeZOhtv0RVZ0xJxVh0
LuJtfTpwS93E8o4oAgY63ENEB++fYtvDgEWLLeQiuX+7uaI2Tfdn1qdm3nb7AzfQzQsefN+ImxPS
Ok7LUOnrKNqJef1upME6DwRM7/ZGOcLKfwC1WkyLcpFaHI8usyNfboSuG9DsJB9jwXRJAnd/kUHt
Df/O/nVNEmaIq5BTfmCq8Tz1j3vLILKzxYcDUarwn4d/5UogbjVWogstpzsoH3uYa+ghBuBXpI8o
sQ/kAuwE64ZbIYPSb7XYpIjf5qXumIkdOJHjivmOXSUmB3XL53mNIjKcf1SA6Jzih6/Rj5t7DPyn
FXywaLWTM5yNsMboTOi41kXNS6dgDo7tsLn7NXJjzLSrGruD3Qs5uMzjV/sLpxWQzcQ+vibtR/Kx
bpKMfaXwr7RzYSV12AV+EybW0jOrEdKPU/bx5txWm7hWoNpZvO6zxFRC3sWe9lymmCQLiqQ66nEr
Mitd2jDYEgxZLrjGVJ0fQ89ns6TH+AyIvAwPbWg4oMnBNm7/jt7dhXkHin1s+daZvd0nvfnFj+ur
3pVGS2gnL2lKN5PlzHkVbFPlA1SHm0q3EbHPMDudDN2CF0J4cXgvamua8Lq3gQZHOuxWjE+c4XgS
5yAMV0MJs/EqEhsPHhhlRuAn8DmbfO2cCvrANYOuPnHvQd86ImFMYhHhSacqS/VMx/Lg85jxn/m4
DGd1fyaQRKozRaPvSwEnsXFjzd+jmcziwRLqEaLU0R9fserPIMxMH+NFNRJN/msZ8zHdZEiCyeCM
bKR8YS+YSoeDN+bIoQ3kd7MZFd+bgkA2fTju1DLsyA7NzZn38URyC1lPBjVaCF5mvzF83KLlHPAv
40rOI64CpKd/9X6ayLqjVdGbdOBKNlxEIg+IWbaHPpdFkjsEi/I5GuZxmDi6+s7G5p7FCAEcXcnz
0lR0oPEci6Mb8vi5+8HWvmRd7ZIg1YcXCU4DSDK7aK9O7qy9a+sIYWPuIU+fAfh4f8mFK8p1Xo/r
aWwtBzMwfnEHFlVXTAute33JWVmG+EvTj7OkJynh4NTGwLOrqIflMefxit5RYVVmSHE8m6/sDLur
nh/hYDyM+qtyfJzV4p3dWuhnt0ae2toSsR+SuUCojnu3cGfCQnqHIwvIvAjvnHz+txFPRfaYQwN6
BhfuTjpcDyPZUheyvgOSZ0YrxSbCnuYirN1GGhnl/k7it404PFfBAXN7rqd2t6jCX/SuevcsDeZZ
BNYb7EB7DxN1PBmXNtaGmYH5GsA5IWzCuIwdqZaD8g3wTOFANIM6idHtYr8iu8+ML5UoDRk08TWT
N54ozvOr6M7tHAQ3dK1mIew9Qsr+yzT8/B0shvcgwHLvAODiOQG+dN3KQvTA2PKD3L7nGzLY3fbp
0PxqBwqfz9GTIJ3BXr0YKln2e2yT/y4ABEVyVtvEYdtXLYfG+Dsjo1CwR8Iak1s9Bo09LIVqRwTG
RK4YHwIKLXhG0tkx1l00vkI5xjbMF8UWPtFd52k3wMvljCqFoUzthbPP5u6bZ6KIdtg38LegsO6U
vDe2QZJ+fO8rPcQaRIHenYENY7G3HFhfyTHuel/FyhDoMU3g4Tv97heAs696APv/DfnfgPDQPVsD
zxqrhjtBpSfZxaGd0fhRlY87Bz9mrw7/HHul3kuA7XgHC7qV0ieVtYgBxXf5vQNgDNRfyjYV7c81
VuQpMkJ8+OnoV4dQGkApu3RKS86auhG+4m1uXJ7WBVd8EsDTltlvhPe84vja4RhJvZUCgRix8Frg
wqHS1VpCsMah1MvDQHECkidtGVdOF40faznUTk0EJLGD2Z4vsnnCSex7dTP1e0ybzk/a1ZbRkpuN
nF/MY6SmkJCW0LZvuZWZqxyvqILCBuRSfVgv6o2iZv9XLvRITQoO24EkFz4iucUr82rtpIaW6l38
UKubkvyaw1WdbG7UgswZWddMiwaKuZGvbF08oLzuDNdLTimpqtPmxpR4v3vILSVsuWDJvZi3yPuq
w13ZK9ME/1jy9Z4y/wF0ALZAz3846cXsHZ0RfGqyIE9oMB+Uu5haWLevYlgI/7ivmaM9GUEcisjq
DcMoKRmz0ldRvAa3BJ/QWw1j7+JgUcIhCrFrVBmt9AL60n37i7W07mBCT97+yT1vZfwMemCbzpfr
46ZDdHhImgJMmmGRccihxkhYfN1WMX3VXiHZMNkpNbOrhlwKe/DghAbV4uUZ2w82VCBy+bHXhDqf
dnJHr6L05juy+3PU/Avj1ZBzk9+mNijUA70BLndZInDYO3NI8WnzhbDX9Ru8VSoT0E36Fqk9nRXt
YFg2Xv1KgNQ//K6zMh+Zff0Y8Ej1vIgW7aL6FlLvI4/YdFd52R0oeWjTIFFhicQkOVD7AAmvEk5g
tEUwgOM2U6yo78C9ZRArjQKuDZUTqQIsulJdLBH9J4qozlkIDbluOHFClgev9pbdQWuQQvcrz7VR
6Zznn2Q7DHRWBRdKCn4aqTWyfh14ssmUIMjyYTPJGuvlEQIIFX0q5dnMt2oOQmqn1x/P9Ga2ZUeP
RafwwuxyRvjczkPHPo240Llqfr8zaZHaSNQdoQ7+KAJ9E2sYNbJ5xsNGyO+fEXPByhSC/lpguUpt
XufgcRdM1xLj/ImFJzHsG2mHQq0UdtHSueYvi/5x0oyJ539fKkiyKH7+OfIj0sejwUYB3aafnTVa
rrlvHQ03WR01PWjo7KmZmJq+WLUKdlJVeaDqFwMYuUY+31rtIN41KB1NIkYsIg2XJYCWkIs2NWFZ
z60wMAJ3RPYnIVkLmHTtI8DsA2aIIBLPf6ydcIl1wKQa4iDGL6fVUv2A4srMMiPPodxQ7h/2zAQu
IcgIj4yrzUJO50skbcZ8u3J333Pmy2v2Er9Heuiwql5ECuFdqX30r2JPb0XtWN5TORlLY6UPAx97
3EAuYKdhyIYm0I8jA05Rz4Ju4R6sRI+N8AVcby/8w5xBOQ3SFmu1i20jx46YiaHUfiBzPBgFljWg
7PTRfeZm80RhHiO417mMK6+ZesZKFwn9rYumnHWmwZjyzMx1b76ZgEb609T7JTxajgIWesv9zF8h
uGXW2j2kYn0QxVj0UjbUgLsOwwAGvV/tsue1rs0mzVlvdJLwwEP0KkDFQEDa6/0BtqE75QP+ymIJ
Z53dlXbHSFb4O+c8Ty3+rh2UqXg3LMWhFsF9qGZyDUr88VYS5BP0mOcaRtPvlIHBNEeQOKazJGYS
jDsaTD04Y4eB/BIE14Cynd96HHu3xJcApB76CtmnVTrJdwOT18qzEKnOrVRrRcbmHFcmfRuFYbta
uqbv1H/10MTIp9phbvw/hp4CjO7QHwMRmdKNfDp5m3fyl9rYcBXemRmdpGvBkodeq9R+8Ota9M9/
rtt6MlbVydL5kcHAKk3R33fluwgPri7JZ/arj3GVtWHI/hExJn0C6wenEwV0wNe7sdYczjKGf3cd
Pogz4ixFWfHA+NC0QPCpI9skSwdCCw9gm0QlU5jEi33epwxLTrjkPIoh8M4HVXf0HBtJx2Rc7QyO
eDoGfRBk9jCguosxaMQr37roRfZ9k/MljkWDP48gEp2r8ebqGFf/vK4j85YT1QYlNyy7AKUnc+s/
PpgtQqSfcEn180y+QVqybqFtoTfblsk5qGT8kJFLdBTWq5THmLu6SG3RwemLtKdtKcLI0j+8RnCX
i+HmxbF5cKGAViqprEJHFCx9UxXsRI7CTj1AARhBMt5EKie2N1McmDmAmX+HvvJr5jqJ4BGwlTCZ
xZMqqx2/27FQmS17Bu+4qHnMTlYCDO1yIF5P5W3WjN+ryq9pKz3qszUadOSs61p3dJ/DkS3upTLT
jfvMsh4tqAifkD/fM0h5DLnjIfw7zDm91GOwlmqZ6QkCvoxruclsYf/qSsyC+2KvpjBTXfBwpJux
wm/g05CWsw26oTw62BqwklgB+UsHj/HEPLYlCE3/Wqoqi5qFNm2x8QVcZcX9yXfabopt3Cde2F6N
CCukiQJ+02beNiNaUrnkvQb2aykM0jtbKj3IZyRYWrew/8VhArwusMPlM5/I/9NnW4MlfbIsaE6K
jJMq5dZ2Amfsavk76Ym2FzB4beyStwc5fXXFy9obDQN1yQhou2wvS7qbH1TPcwoXEUgPm3iA5i24
tc0QlMZpbyojbHJjmNYsNCNCN2MebVH4bbsK+H20Tm74QhqtAHsKTSzAoHUW9ksfHrgu2+5CalX1
j87c5jxZqtNM/noG8U2IZqjXUEfx0TzlFQP8Qg6LUH7TWZgA1H8+HtG/0cptD7yFXG22/iC5Xyc1
FGMxesVEZeeXe94LbbCREKyOWT5Bgij8OUtI0A4HXv0jznTMM9hhzp+eeDE6q5vJMWbtRTjLCkEq
Mhd4MeDaeeumnpe57evxk+xZUmYuJhtbPP/p8prDKJygQL07cOhTCwpix6+Wj3oKHXJBduAIBNTT
zNcwHlIgobeefOKPtxEAJqRidbwnnXxS+kB0gQSJiq87dOxZB6RjlSxeWPGELNAifo+8ERuqmNM+
ctdHrZmWeeCSfgSdQTMH9PXRNbAocFo8hJs0XD4NA+0CoD+O2eLNl/hN5xBsCghEirC5FwB7GcfY
uriZuOvjXO5OIwTH2xfNIv6zmPNKnansDddQyeaJk/6Qmrsw/4QdA3IdnAtYMqLzEBn2JZoYvkCr
vPeSQ8lEYm+SsWreFr7bTOwVBRC+lw77YH7NOujxiW76K1eFmli66Nc7xS3YvXZo7exoaGoF7QaC
+Jttn4zNN07w3hQ08jUeWp9KT1RroupeLeSD+2R2RmpQ3H7ma7luqr1uhHkcox4+urnmQ4etg7H0
nERelhDXLs/nv4KuRJXHCMu3EiiOW7lnXApjv8e0n7Iuv5bc8K0jm6a+sJvnjxrZUxOWULmFixpa
GxvyfDRy5sNnGiKmrz2YSTjD63XVoxRU7wEydRa/BpUEX3BFTlkgKxc/xQ+O7fcREt0WyC9Ncv0h
XfcYG0h/RGLz6kVI4tRBEKSds7mCSG1SEM2p7rGbkcLsJBAhPTokEKreuxRxoZWPvpFK9r9VjDkk
ibsLpuFz7XmbuBXE97v1t8gyI0JLdegf36K+Lm4SuGMenEi4Z3lP6enhh0/dsAPsV8Yrbv4GGc0E
JC+jKWqxnzspuxJZzQKngFkUxcj69nj/01XPVpYvPZk1lwgH0aQgnD1MCTKA7hcpCP5W47LG9D6R
snN51rvP+T6GIwpfHqpaiOBzbZ8wsQMrtsXSD5JXaOW+xSPIWi9TTIYwaWW/nzZuKegmvvDVdYm7
7aN0y1EFiJNkIeXtZwABcW1f6g7B9n82910JD4d8NPm8fLELxQpOJjVt8ctE6R5WUL2t/aSwLA2f
x3THTqXZk4fAr3PyRwJVZ/VYrdLautQ+3aYP2uLctTOuWeJzCauxQ0yW5LzRhPY/mEmbzlxo9dbe
RdljHBYuGzmz++DLbpoc3yLu9e6w7GXvawjqYfTpFaUxD0u8cduarGY5HJJBg+rCo0Hc3LMcknMo
TfiobasOLyiEpEES4E8yWBsk+4M3uDNuHbXS+RmB+BeFa7eHypnDW11uhl0KFTmJN5xkuuzcVmUB
ZJprw8pUSbLwiAuKF0/oxAMTVRktzuxM/t3kmKY6XiFSrx24XQKEqqtIVvY3FKO2LfnA2pNIhjKG
1s6c7p8EvjREOhonkut+tPjLtkEdroVHACMjgGTehhg6S+QcPCJb54td4KHQFfe6ERZcV6nI7yaP
jBg7mTPUiKEWek5G3Za7CKgh1AmHzD5c1vPZp7pg1KOomw3Kq/9odz7qzXdeb5yKqqLS+cMXJ8VG
BYcAiUaClrXhI+fjk+SiukoFVLVg96Yca81lGBED467+94fBWhL4HN7Kqr1KkhnLqtS6XfhM66af
dVqKSM25GT+88dqRMyHTpV+pm04kXnSShbYulQvprhsnm4KKJ6UzcBetQmy6XZkzSv30xMUKuOvQ
ty02xTCHiHYlf9YRXahj2etXse2dxpwyEkOVciMB7pagWP/phHFlHzcMvhK3GIIYh132KmGkxBKg
gDXOC8F+xRrr7sPgqEAAjZsftj5VasOu9fDTxQ66exA1q6y2GgfPGJV9fsDIV9ETmnSjUrNWuafB
7MH355uaEG/7zE3iyt6s5Db5hjQg6TUTBwI+XFCvR9lW539B0nA+kWXYXmXDzBSSo9Vink/URNvA
HrxghybxCY9gH/VKHB87oHL9erFxND57gTXz+9u+2ARvRj8Fv9wMULayEapHDdKFHHX2pwMOoiSv
mlq2R1ruxpPBv98iso694YCpd/hfkx+VGjrRk5Zuvs26n4jkZ7V2TPK2QuFKuJUazupndtx9U1q6
YhKk3CVCM/NQq23mek0aWa0TA/jkFmLMQMI0llsJm/JxNklUMB/WlHDqQGIYiZE8GcDJdFA9pkl4
G8nhFsiboZm4jHFRGGMYPRnnK3BlMoecARDIaC9NS5eiH/etC30DEoY6DzpRhLfBp8vSJ27/G84D
P3xSWvqC3fbiH1kXqSlRTVfu0xonHKKSRFfFi2Llkl1XuNSS2nRjkxLD7ZH3aeQ/gosHgDUAyQn+
PETJ38cqi666OHoUGgpjgRmmN81+lJ7j/7IyNfezrYWPP8DvQSafgpAdkyj+60Rjyfvi/8e+o+ts
J6+3o7TMrY1MlBWGzCVIP4mq6c8uoLFBaYh8eUDs/Fd/RVFGI0mx5o4+IQWnXwHXPefu4NhRzSa9
Ikly30Tjb+VuqJ1uyvj/LM7qb0U5BdM2aC6wr19SiU6hkpoFiWDb7kX9DB6nCApNDatFClg5vJps
HWetKjLXcTG59N8eKjUGnossIiuXbI83qgdOBsIsy0axBvzI4NMrJVTYyNLrC6BqrK/VJ2/duEnR
/aNP7cnF1cWiLTrabpC+HtcADYBhDuO50x8LP6EGP7saaHyWaatqphBIl5dVfiX1VkL1YMGvGfRc
NoN7/sO9kwRek1Q1YMJcsXTLnlfEU78TJc1eudqe7crJrsqS4S/khhlicS86k7LEQznTiytiIA76
rKxMtfJ6DC2xeWnV0rIPlpHdF4DEtLajhJkoFeam39bdsj1oiptu4WfUh0hXJy1cgy1VUc6Z8WY4
7j79M7uJqS+USsoYft64z0hsEjOgDaJo7Zz2wgrdbcdenu//t2E1Tm3uCYYkSnuLYK4gYzz6MmCT
A3lRAMHMQHWJmlwu9kBVjYqj/XKon3PGHTNfHHByk4enoOi1pUF6i6AuX8x/LNLDohkZDE0yXXTj
YipK4yF2CrAVdKR6odw5sxJwf970O54MsZuBG+3PcTn6+h16dn0FugWzKS9VCmhsR1Dt0oq7oVhW
n59D7k/S0jujZ/hbO/U47VBTdgOy+PVTuYFie/vWL+O8vKiWVMMojP1T1rlJlGr4THVPFGjyrRIv
AuoIPz+u4neaY3CdyYcJrQ6BxIRogtIhpeTgs1tvEcKCQaoAddD8PyTjwnc1GFSXcZ7ijYrbQpjm
AnvlBgOmmDKiqG440osKhwdJeKcmqWxkYCDRGkmYcyS4rgMVCshCHjjH4vQY8ymgKKNkehzZA8P9
NXHhzlayRpogzsK48N8d42qOkHZ6tu4Mi9z3n4UzcgdGJOsLUpnGFgYRs6AgBaw4U7dzRQZKCpoR
5h9rt4JNkjycj4FYUCykXJ34cQ5cMQeZrFpiPlmvhqPT+UNy67ltNfkVq8j9I03QQXbZq5cM7Dpo
gBnQ+W5Yqvu7PwO0d5IJ+deb/Jj7Kbm4/NCB1Px1RwfoZH2bZPtP5Zog7O2DF5VUJsR1JeEmEaKH
qSVZddXHyFIvsHYOO7e+UcHlJNAEXs8BjJR3eNI6Tyaa1uY9Qb23hU60yYCQ6Lmxj8FwMhWQpV6P
sGr3M+EMN8HkwIEJReM+rkUuhLutMWbzhEsE+yRRwWOKKseApL9fXKJ3OYnUCo6hv8J/H7/gUA2t
GsYjLt6vTNWVafrkkgrwJMIv3wkhFibVjkPGh8FVcmtLYFKST2cRcvGrYlObYxsX9onDJWi/AkzW
OUYjxwJgNSM5xLdqNdB6+4pGWdlv436ormOTkT8fzxzaU9KGQWwRRGQrC5r2R6i0OBptzoP3mkr+
O8j4dq3Hc7Vb7cEZd3Tx/9QraEdm83xTvt0aY50aJ8wfdTBJglLC49GqFm3mV+jpZ4RwjrAQ4XJa
Qhpz8IH8+vRDQK7RKzzOeFQJctQHZ6IKFPxfih2rg3lQGaOcP+caFEZfHlcTfD3GR5F2r4HUsesv
D9C3VGYjQqhWaqw54HZ0VeyxiMybRMLMzcSngFEut2mo6JY25rAZ3UbS6UsfVgl68sx6pbH/VXJo
gjlUUCsOGluqlkj6ycdbET0pRR3oyD2EObXEfKG/AyHIs/W7OksGreHaFk/oTCpUu1b36/qAeDOo
5Mnppyji+7R0NUMH3fa5fpy7JlFV+Lsu11QwR2kt9aIljtN/o0iU93XXbFLdmPhUOWDpa+PL7yik
q0tPBcFsgxoJJPZjhM3FbSK5Zf8lGEGpIrwRrggufuGw16D5qwB9pZdYUC7mCelgFj3OSC9L4CtW
F6a4n3iL6/jvhZf000dYDrReHK6clbbVJOjk9e9wgHI3mDzzX2dOTka3zxnZr8W3akNjj9uwUqSX
GrnltZOafn9ruS7cjhmU/lBqMumgr5BR0c2o9YWOND12ZyxcMyLpcIGAdMPozZfd9aEZkdVChmz9
OgAd73Qf7RAFVJ0UMHEAGSXVCseSYKWREktAKoL8Rpjf48Eut15eN8X5EojEJuBr26lSjOSSakvz
+hGJoiJ//CnIJWmv9Ha4DSnsYWA6HFo8tHdE3fhBy81bzRlniOGMdKHgOp8TafykCJOMweQ96CIr
13VDljjrsNR+IU8Ihfa/whWwwOSeHMjiWQf1UWEjpw0/Th1dWXFjN92sw7udvnsQw39KqeRPZ6LM
v2Q7oT+9JMW2avsHgsz9xWPTgvh08PnToElp8hvjoneOQRnSds8T5kTuKBkxPJpA4ozpQhiluB+T
CvBpsPtvih3+d5AWRodnqjEoU4zVixdl8/7vqkDCFbQexQGIjzVaHvyLYHHKY/8DWQpj9L4RYtGa
AhhwKJvAaPBXKRHwEvljj4DwXUDbqN1Fp1qnTLT/TZ2X15SfWC0RWGqqaG5dzyIW/9VHsMcXixJv
j2Ve0L4GdzTloMG5MyiYlKpgeqr+kVJ70goUAb1YHfihtuByrS24buwik6sx90GjlgeV7TRUgYe6
F5a5fslF8QhE9hMcRLCFOGC/NMiLcrXtjUA0IcwTU+9PEO/gpw2G5saWT2Ue0uCQf5ydr1Kh9QSA
Om5OZaJKtubwVz9rxeuoINt0MKQp5zt+jnYxqG0q3WqUPy3jSBY6rso7+x96SAuNYyn6Lmyi8iCD
CzdGVtiP9sQinWN37dBGallN8yQmxQTJQqOTCTyyH4Ry6OC8ZA4YVEzYdIY2oo5E9HOqlzsnsh+2
F/keDKDLX2ExWx8Zi24wAfKeSUd2S/GpOdjvLCoVDC+NJ39y6RSft2ChXgPzBg9rnviXu2gOCmqZ
qs3cgqv+sVjn7jCS2jsKBkFwVfOMTDeS6BXCUAxscdCdsJey4lbbDMzQK2S4ulbqSIeZo+B15RzU
mCIo8qn1UXWdrgKKdqq0Z7lt7i1DtArg5sBXflA3ukGl+DSiQtBO+MJgIJRjt9T6XBeBal12Ijsj
NU+UTRoSjfQcM5FTCTrMpq4zN4AhT55Q5sTSpYYQF4f7PgPVdREopqHaWKjKF5b8EmPBiCwQpDZ1
+E4ocZ7F84akYdlB7qXAdU5JhCviYeEgLg7ZFFKdXRNtXCguLjbZd2mUmoW/4atcV4L17c2JxItC
7LEVSr7otYkYVMISBQB0lw0LOMHMj+eok9RhenWCetNdN3/SRolmokAsOsZ+K7Zp4aD87J8yXfeV
XYSHXi/mcn202XqppcNrqrQQ/HRtIA2u1S8Tzs+9G/7LOkbo3mh+mgAOixYM5UHDvdf/OPwln6dy
5NXIeAUkSbYIOzZYcC3Q9DF4MK/0VgUoNuUe9dK6ughHCcDEpO5L4GWWM4cU16Jayl4m1fqLUskD
P19X3Gj8c+O0QhzgZEowRJj4urMrKNMcQYoUBIRQ5f06XHQwW00d5NlTAafwrrGj1X/X+EEw1FBp
9kSqrsxT7kiB9t+MaTF2D5K0lkZF3K5bo5pvit10p/MFhvJcik5SA0oS9sXzJjE+YkQVWpptphXs
OQ6VAUWW/C+tHcDN752x8i/GmEbsSN4TDgtWyiidUX8DD+cuO+k2CKIUVKKCzrzrHrXr/pK/Jt7Z
+mErfMsNiQrn+Mg+sU4gr8uai6OJatCMdVdS6L4nmVDyckwWgkE2/Fn4Ald0ytn4oBXVO+qU0jAh
ru0/fxHU/1n6B/jgUytiRrYoywUSv3wUuKnrDotn/fkkCbwYIlFwpEBp2qgn/KXpduIBHWUSqEGp
6WSTrmV1KQmYzrqsqBy57MGE+Jsvt8RubaVZRb8U57BAagA2UolFmJlZn9fhEy0FjcBLkk7zEOE3
5nqsNCUABkYEgAYwQpRB+ZS0CoyxB9PeO3T7kce+wU6rXh4cAuof/j48fOdRD8lWMaxtkENh2qkc
SUKAgvj5MLWJOn1DQJlhUpGaVoCM5JzhRoKh89UZacS0Rylv6TCRmAlNwFigeVJ8hmzuRMp7ckwf
OoWhr66xFkMqPHbxDzMMXbioiJUXvk7z7h1cemv6FarZd0hsQnv1SmUDe2/qsqBjv/Ewvr4yxId0
dfnpi2KqGAcygpAKaISX3y35q+xBp+xKo1FOk0ASh7LK+NOcQs/rBMzqZdhd03WRJS/uvERaF6Qi
BsFTMbyom07p2ffuzP8sjU3T2O0khlFtkAW9+H0C22BaIgcvmDIULk8vw2CGrR5yW1cnRtec1feu
TYFbfj8AlPjhO9oT8voUb6feQc0I+LTZ6A189Km/sFycs6bBk0qpz61MnrbD6hdmRE/XY214wFeQ
fS+ZcAGYgxHOcItenzAC52loWGp/5+RFzT2hUwvAEqo2fSfGMBWQupt6gGfSXc2pjf18N8FpdsXA
92pK/I8h7ndWVRAnstfc0XcVUuYkp12aWJNJ4GYDeCwwFVBvk7Pet6UMrEF/8UGMJ8/JijT36kQZ
0SLS6llCOkCwQ4ZDV9u1fHwsA+6Egm6xSVyzFj/w8j+Uuu2sotSp4cFy6GQeZQw0hB/yDoWJwmFH
wpgGOAhyZoNGdgArTGuIVpaQrG6sH3f9O67JxmoB23m73xhck1GslAGhklsVWh1SHsEQw7m/i1Qe
Ii4scqS2fJzyrjzgCD/kKuQYzS6v+M8ZuDcd4sj+3Dc5SII/jXnMG/E/9pxfCvTU5kbgp2TgMnxt
TftwV/baWjc3vEGwgnGBDMKc9NJHvcz9MbLd1lcpHHjxtzj5R9maUHFducJ+KTZ6NTK6HbAtmUyl
Ek+mDHAEx+S+EFuDop6PpnN/c/kNNcNBQ6ekRT5xbXgzHwPnftNw6irSWOAvjPUUEtRxqqi+81GT
i1p7WNY7zQZjkOvALE94BMNuWWW8BuDjSo4K1yEAn8xVPM/04FlIe0vP0JWFSQsYr7g5y7nUBRuj
Ij4ZBXkruYsNcXD4YI3sW/m95Hg8g+GlSzy7jjKsNWgNKJvavYyCLBVyf7FSAZ3JRfh3FSv67TGA
LWaRA0IdZvZeMgS/wgBEyPEar6zf2jyqcfGAEdAwR+crmByPtUEM7F3zhmnyRHfQKF5HVNeb1Kzs
D96Jwxsty/3Qix751bsQ5vEQf2aYV3tITAy05qXAiaqysvQ3Bq5cCUfrrmsq1nq6EjzFR5xe7Ni/
RsN+M5B+Xs4WAjXPzsc6VZm4bMc/VizTs4lnGzfpzBGczN7AmmQVbNJbRHGa2vccaUlAC+VsrBsH
B4AMHNp5YGy8ZfKJu4DmPXS6VIwSIxy1yrgR3F3fKfBjpbNoNBsw3AMyUJirzYC2KKRZ3MbBysmJ
GSf8vHM9Gr0Ba6An3pfgAN7CZ9QnPDjeQeuT1iaPpuVq/OeQXtkXTt7KV1Epi2AvR+0PdBcizo4j
BbnhiDadlo8DvKHgTTs98n7hEWI4BfnF1EPimaB3s3SEMO+9fzKsKLbXzyEpso13EDltYt/sSdFp
zINZn/qWoL+h5di44v7NtNbWKEcImj3kZq6T+yRpmoCTTO+Pqf6G+vTxjIe8IWD77ZXilCMNm3lL
ltNxdhbLwOpTYq+H1NI99InnfTT/ZKH5lDe9jgpjU+axsdVr1e1Y7Gx4tAMC1qZNR2Rqlu21jU0d
WRx/2yoVsBR/inrrnGe44AyoRFhKTRX6qwg/k+tGDjCknsIAg5FTBMEsHXOaQ4O6w7VpbTmS7Rn5
/sDtk7VV//P+Wp0BUYsR2HkIGgh1Wh3oCYavqgvNGrJUfkJtQnhY+rsUYvZfZWmpK+ka1MaKZ002
xQT2mqTBeTbRDGAw3dFLyVMfz51nv0ImYgXPwQ9RdSyiHPpw1WwOAHNY743eTkbDuNJROPJtL/fZ
qAJNpfK2qLWmTQWePC3hTNbqK8XhuWOVIpwHWObxOJDjrJhquYFY/Jf3V6+V62P62xj8SezvNvhB
zCa3TFzHZfcgyV4fzZsvjAquACx63nSYhxV0eyfljUpiqXxDkP384hrlQkLyoVWjTNrGFOW3DBui
RXyM6ssov4OslYyR165NXjcBJ/kJsZAnCioPyM7rSNCyyBniQailmKE/KBLd8ATFGUF1gwtNYFKL
RsxpT7m66HvBTwiBoGVFH/nXxqkfbclv5F7iHxunkIqMz+bWSPj7qyojUwT5uGzWnywnku1yMgFV
SrAxYODKx6EGePgD+SBh2TojGJyzacEsv9J5XaB0rRI+jlKg30lMsE4A2Si8WX1JmhndCfuL9O2R
n4yxr5vWs8C4z9k0MVmzksMUkOP4+N4bR/hLzTTgCm3k6FqI2wJhItHfy0zdejIKf8RetGzooEYS
swF5M1MSgqcRkWBLP8Kh8DkUbHrw1Oa44uJ9MeHCfFeL6OUgnNcVyb6B73aZ4Qb0Fd8Gld1cAC/d
24/VBWtO1QUJakxIi7vxfCXJpM/qvxLdim+YKD51qSGV2nd3Lgrt9ClpltqYXPoAql2VgzEIIMmS
qQOIYTryHXoKfIhdZbVSqYR81dlDFpT0UP9xGvTG6KVgnapHW7JL0EzOQdOQtA0wAYYVRKstyfDw
BvdL1H4YUjEN15IZIM2zaEK0rNLiB+l/7b7eZ320amoJaQcXYAtqRkBO2nIXcMgmFf8FgtoPkX49
pTZhQd9gbrevUMWrB9S1erT3tSJPhQhqK2ksl/y2WUECZTD1z8PILhkO/QS8pdRvcIOxbkTcDht8
9sMgp1cNjTEglT4riOwhhMdq+C368zDswQjvtXCzAbA9e6eoDm09JQ4Qpkt+/7GG/VruwxS5MscI
xP+YBX6Ca+Bl/KXwHKDLYN02NZQcER38EQiyLrjVPMtCnudohoJjC/lzvZaOaN1P1TF7Yzr2RISd
39DlYYolB7LUEKZOnQHAEqhrMgz40vAPsD6nwlFgcNVzXJy38itPJb59BJobtwFRJMC58wf0PjFx
qtbFKAo48wwttDEnA2qKxRrIsTp3ARkwzFkMS81QpOL2SOXqV5UM5e0oq9Rz6WpsIfMndMB8Is28
gdOfP0cOpYGISU8qecvGQNU8KkEqHw1+kOpXFIBv+I0e0kG2DLHz5Dn+hbsTA/9dBpjGtfFpFu+L
/4BlQUGq/PBzK+joh1238GRb8HfHl9QXWWfM71XrKWJmyFYB5WUOCjvqY4jf/kMFgOksTlilMoT0
LFy29VQUE0Q/gIkrLUG0WlmOP0sAo+tXYmpBOzs8Z6yKuZfe+AolMAlKuQLTTEV20VypWrSNOaoj
5aiC0JMBaH58JxPQ1t26VntXHvQpC+j+six+0IDsr4AV6JLcH2uKqnly080qWW1RpuXoOtciuzjH
99gChgSQjl/11HWCikFp9vlO6c+Ch36Bb3lHQHLbrM2rw9FiHKqe3csMA6XvcYtuE0XKOMyJyRRl
TxuiVLbETve6KnFgQB/9somglCnXyGu+q1wsLezAkv7uBLe/2MTjk36GL4YPuqp6C4rkI2DOgCr2
aJEPJJmB/tVDS9YHWn62yREreZLgWZk1sR6SIl2yY3XRtfUzvJOeEHuCx6zO7GV4xC4unPu64C/q
5Xc9yQGXg7hyRrGmFmev+lSjio7UVxNYeaQ2PzZ2Mloz4uEau437qFXmDSCeHo/B+/WStS0Tx44b
iZSvQBOMnh/CD0HefP+RNA76s8hXhK03+ukL4Z1eiKkAbWtSwvVhslrCIjnOkzYY0pfz7YE8cT5O
n8QQLBs+6K1nEESr6iKnhYLSi3Y5CeZpDTZ2GSuIsa+zvARfbKUSb26ypdQskChFqM/EWrfNz3g5
RVA1wlxtTnFn8q4GplMMBUoGcnfL044on5d2aPCov/ol4QtixZMFZ0Xx7//Lgb6acDS07Aya7QtZ
KpxoKvroHudH7AtbVopBuc6JoBxdTbFT5XLNhz/8jn3diL922PQWFNjVwBvGTNZSsGy+1iOGppOL
xo+FnTjbfx42HLph+CkvZoxJ9RgG1uYg9kpYV17YhFGjhlceNHRhvNUGNbczPdHWZGkjvTvLXaYT
p4He1aeJbiPA/AXvQqsD9475Zn6Diq5j0Mv1dRQaytOt0z1myitXGAmR7lTaO2CgqK8SqpSMpGLZ
HRhOpcR+J7MRQjO4DicEQddOzeItdddKDm303wP7PfoMuKrvhJj6IXO5SzP+FCjWYyYreP8phy9r
+gYN2GTfUzQkMjkvVmSJ6LJeu7wMHrqh0e57loaf2urvGASDwnGG2QScrXpoMwEyNvRvowXw914o
0e7LV+0kdVBkaKRjmz+0aA/B7gnQKg68XZDDJcfe7G8xNG6NfHbgSThyjteJmrBQaCXUN5/S9TeX
jfa+wkyBv/u7BiDjALgXY8sr3Q+NHeQCZpy9kVft6RBz5IWMdnxPhjGgJhP1cpthWhHOMr/pbDHy
3uZ6h59YtTCGGYOk5ZHuRxgVSo2TornaiIwcyn4cZS3AL/9fnDY5546B4/Vlf/d9BrHM2vw9jp5A
BlxhOjm06cr2MV5AbFvx8hvkGqY7mPP+0AmuL09wd3vK4Kawf/y1HuztndvqfZhJABYUO/lcwO46
c8aC9dNADkEO6KiB2ab0Y/621Ndh+S8GAeL7qamoV6IUpDJhksFX41KueuqJ2lP/kjwqQ/YaSI7H
Cy76eUyqByg7dKKKGnh8DqQYwRWov08ZuT3ozGHIqHIYykQnh5Nh6uoGQDVfTWlT89s2DT8D3u8A
lhfr2glwoFVRop7s5eo+njJHyqkb/NLuhcfekIThJLCIQ1uJAk4mXIXjdtrmzQyl8tktz4XppyO1
9Rjjsyur4kSxr94Lv2KQAp0EBQ7V+RrGujILFnEa4lLbe4ack0fwbmhchRfRyWfiy0NkdPuKs9AF
QhRf/JpHSKXZav7x1x3/DZInm4eOtCHwCiUwRSd/UB93HWvoc90Q7iyzfagI8P2hjlLT2bUQexN0
DiENHnxdLbUOq+8G8q0nTFi3UH6DmODvtsKO93vx73lzocJ4aD7q46oKjDe3myhdKVmBnY4HglaR
V7mr5tA4Y1YAHGtNOcqVAFmZw9FQACIp6lPK2294IJ0kegJd5OYVdKkwwXOo+qF+Vbxd3wOpvAQT
saF73Io4kcnW3uD+RPbQv3+1kr88NJKk6S3vxpCDp+KLRriAQxjbEWy8oj9PLs1bgdLP4c1pAGSk
pXYhfeKqlAvDok7NmCuKkDSjAIVwHWt+Pexg22YpdtLrWSFS3K+axfQM99WXbT7m1o+Q08//iLb/
AYwfW12G4Hz7Ox2vMfhMioJWw9f9fGNDzEqsD3SMEpzopXX+UzMExwaSCfvTDntL2LWDaMVVC8rJ
6fMgEREWjtJ2QD87FChDKqSh82CRULMHljXpjC4Y3Hiv3b0xDKji2+uXychZ5NPmY3CzymTt0b0p
uXOz2A8SsQBvSvzdZI8r7XuJ0tMq8QKE5IFJDYrc7g+K0WAAxUutHb4vc83DM5SVnWPf9S//j5Xg
+5fpDZBI4P71r5ESyjXGn4eb0u63ecxATaqgKkLZ+kIZmsbgyFpvq4Sf9zZm6gGJdT5tChKTsZol
p8uLzgydIVob7MCLXy7pTsqvJoJIyUXaFLYIoyyIUHQhQBQ4mtfJfeRC9j/slJfyuwMs4bpZtiaI
oeBpJQmz4nn9Re1oHLJkZ+cJo6Q/pBArNxngeclOijWBGbH9S1/6WO35BF1I0mMgbPQIJWgrYzfP
Cp19HBwpzQfFHBVWSczfzs0gp3ktiLQ08NebjZB7TbcUHKEh/bOvQPjLlBfeSlAvMkKmHB5U8LX8
KgdRz4SoDTuFaQjCD0aqUPB6LcMCikWaqSj9PZkyq1USs8wugbK9cWSchAbAweJa4C86Dan/Wr6X
YvICSGPL9gXQ/RIQTcZ9rLU/wr2ILgkbP9zpQ0cqtviteFu87k6yzTBB59xBRlXf0lxO8HLVu602
0P81GcoerfYJ/7uH5ZjNeZ6A6r9gx3kc3Q7jmkR/NDuhik6bCJxPLElVXFQkHxmGaSQJOqzgiNjR
wgCx2ogn4qPsYGqeVrmF2+2Di1TpQoXXFp57+hWOJhYzCz2M15J7ElC6S1dPFg+umzMotda46rQe
cCFdV4BzS9+7U+UU2XNr2Qfb0DLmVvKvZ4/UMTaMAIsmKWyQrTYGQh4jj0FF/n4kd+5+slnAKEPa
N3oAFbuBs65/WqlbUwJmsUrrsg6H8KLi+dvTXVNqfH8c3P5Nivjs8R+jwLB1eN5jyGi40Eax08wI
ppMVNnGYEx/A4Fqj8a5Vi/L3M7QBb6K60sJADvfSiCY6AE502TRVMpr9+7JjnwmBK12kEUZEzW7W
uNiitScu0DWmDDbmyFudG8cv+cygqgEcn8q/MSX+qTolfts8pqQoZYAcCL63pG0v4Uynm6MKWACn
fYUzFV1Zr+ATCKXcUGK9DJR5PF+0xCSAWcsQk6PQQ/3p/uagTVolVQho7Z4Vq9KPrA+BrXnE7hG1
iOpDgzztcChqgWztL+UauJcevRdri7DZ3dl1zyGuLBCF90NNwRnxkRryCFNN+0S0MHhIPe1ZD1lV
TUj3uFZEQJAjeXvXv7xtYWaf52pgy2I5VSnEkINWRnqnADFH6OT+toeepe543toXPknsGEiZrlBX
d+eNMNzSNFKKUC/eFMsA7GBh1ibrw3B0LgeDg2VJQJxW3fGB7ZCqA50I8d7WyPw1CctAPlyWiaRk
lFJiZw7+cN7Q0GMYyEmE4b4nPD+Rt79z/q6Fxi/nl+rcsyjtb3S+U4lD3qVxNzacWPNAB3hvYRlw
DfCoxI1RvroKemzbOJTjP6DMMovFLq61S0artIpQEGSk9WifGVV64JwJn7Qf3JkV00kWZFfbb2b+
fuN7S4XAEDubu2WAstdUg695gMPtGV0eZ5mdxHgGkEcQ/FDeLwFZuBpoMR05KOXxjZqrPuJG7q6k
590ahpEfpfkEJmfjQibocAujdV2yrm4yNGn/9yqFuguEdx7VDjEF+4INSmVjRxa7EdyreeNhvPoS
AnPynG+cMEflmh4uvDhYwzu7QrBSxBVBvM9NJVwP3u17+XOoGJLxPeR58VN2xU3GEIGJv/nO8Dmf
a0Ym24Og8sgyAiBak4Yr3XjIeWVdEgQn0qAqph+QeUlP47g0/qc/Pw8rRaQWcI/fTixm852dR7iw
FKMrCHBRHTk+0StCwObmDwWneXj0fBuMtV5STK0OsHAgblOz3zS43nmRe590NdtQsgJ30IWcrC4g
4cqsiKU6Mu5G/d6JWyswjqq0Hx9hj+CH1BHgG8rgixc1dB/seB3VyVdRWf/BedTFdHVdwDPozahP
mreMe1YoVFnoNsLkd+IdDMhYoB2j6XEoVYDxM9gPc/7/SI4Z4A0WuIcHPGHWipwXnvpNRnWlgG6b
mvNTvrGWz1yso+WzG9hQmZvaipK8XZWIlMWgurzWYVx/5MXgUdLD0nLO/XJFstHrsC01QDuH7Vo/
qe8p4PZFOdig2+ap/sNfEASuxKZwnC3EinSrIktMw2E0ofTfYwo32OjImSoRltFbcehwji54uJWO
EEYbYNjbSqEyfdVmi8xzKaTJAOG5AgvEn4WwP8J28I9DliY4UEYPHKzFSNps5DJC8AcZYd7N4UXf
Yf3cDGPtBZTy1t43a71FmLhmSkFij4nf7yrg78PRzGPqOErEEtLRyyj/fwvTzq1DQm+tqWOfhk6y
f99HbNmueWda1Y5WzuB9/XCSlWdRwgIMsMkdoTQV0K7hs1uAPjtNS7kUfEIGahOUlJJrw9DY0HHP
O4wEjVDFc20qiDY+O4vBTRwv7xabkDfGeCzqPHYJDlFsAY9MGzSwcZBeEmFO+1igoYH1DVa5VigT
XpE0XnJN02P7+HAOODlGF5dJbWpTz6vL3wTqRJW4u2WiUkc6ktTbmxVVzNXh3CMUvLd7nhMO5+Os
xU34ZbQf1WhfFvUxZ54pfY4kBqodkvRBC2iyl805je2hBuH4CNxyu1AmlT7K4Pm2w0S1XqRGhaao
47fhQsZ4+kKRyLj+z6NF+jX3upWQ1cIeVkgfGvOBa09fmSlri+mPySlYUhp9Q+O/70xYkXzLnSzr
zObUqe1e5k3eRGRvIdiB1l8Fxdj9w/k2kVw0jMOmSSVay1LmOYPrn7E7IV49TQgGJOiUpUBtSYzj
I219djdZWgSfqHlx0WyLBU/23P+Z4dfNz0vN7tmGsahcZFhCulIi1Z2JmObKoAmZr4ie9ghK9DnE
nrGq/DeKCj39yZUPMwacRH3aukCScg81nd6HY9CqK0WQfWLC7/uiUpkbDm5wcMZIsLnFcGJ3PeCY
0xEnKOfgbqXFAXoFAR+BXD/+iGw0ANX2TUm0gyU5jbnpMDJSIzWa+4bg8vrs9aE8BxURu5yIoITS
OQ0gRIhGhrdb7S88m+vK/oY3Fn/EHQb+EW684qCt71fZrdBW5DDXIb5CE0rpGtYQOfLVXATkTdie
KMJr/h1qjqQ06850SH1Yy9QcWjO97k5nmZTnj1chym73GCPJrqMQUp9SprRSH2U/c1PyR5RHmctQ
JjOawMiZyQ1m6bVTN3bVth44DI+btcckxZY3HrQsQkR/PGfDbWPYio/c/EcAPiMJWIeYpNgerBi+
vRM5yP2PHCBLl09mlfOnNJ6FHevoVArneL1ce0cegA7lzoMWjxBndfSiBFbSNv0zLLGO53JU0sWs
Md3ftNDY6eu51MsEJfMNJKCFfCdqGXW/B4FtMZRXmXz41BC4ZtBNDouC9f2Ykx5LbRZcNGpvBAdu
o8b1nzIm14mwKJlpn2jUw+uBuHi4IJ7UVECXSc9xNe3uO5URC01OlGa634ndnS23cYPF0jvwdjjW
PKnUxS53mvUULmCDlnmvSOy5SfQ/eCpAG5tKGbeWvj3AD6yKrchpk/SWe5DUi7vQ4m5Xk0xODLV+
Y6LUigDRa3zwPBCyJuydjdvRc9OdeIzCiz3lQ4JyyPJ7NgzOjAbh3Zp1njKgsZIqXrIeJ8+TlkJ0
D9B4pOWyQU+ZxofjkdDGq8vFJ1TUdF2hv95r77qmsAmVhUNbq8fLZf7+Evf4IvOWOxCfgR4bjvqj
CPP7mjPR6ASMbFlpQi2QVdVD07dLENsmnlOMPhryE9plXMoJcZxw63eBOcMhN2v4oQzS4Uq35Xqp
xnVy4ucMknInscKLU9M926M9Lx8ygzHTu2Q/OOOd2h0TGmDrf2CavcQVEw/ij2TEvrbN89ezTY8F
jrVXyH9kobc6ZWAGVUnnho/KHufs7kGxlegg8AVcV5h4RZbekizcW3p/qeBnel39ZlousyL3qUUj
6sGOaXFZu+rjTkORNrm4UlSELxw82bXfGvpCuDoXI+JvUtES9pBTlbDibpJ1p02UDTTDXJxp9vxF
L7/aMB2SaqaciPFOgM/gaOZMG6ygrecppA/NsZeXRJkPfhfPtteNmCfWGz3bTkDI6jaJKeRPHcId
TOIPxihm62ngAiD8rCCrE9Flwk8hizOCfikTnVt/pfx+/MeCxpNm08mgwe0XQcrJoGVKfWeyhCgK
knfAxRSd5SoESScGBa9JCQ/AWZcgbTQNlTr5UxneoWZaQeVgak9nnNQ2Y9Nf44zVQzvcPbll/w3i
tEL4l/4WMERt7l95TPz8dtOUaEtQa5fxQn0NUXRm21WLs9SdfQ9W7aUp65vgfdyb/xjV2DxoM8BI
PGu69yT+fzeOSdJpXZJqbGSaZQImNrfg4ieXxRKand5FG8ePkniTXlm5zmdyA88kMMELRoIL5ZOv
hia22zCPHr7BW1PnwBVdhoaHZjWNugCXxxx4nUWdY2yqTqEVZ3MaMhcwDeZtENSfdYbYz5PPgast
UVNbDXawsAuO0/Orv4hBmghOB/OZAP2WhfyQfBnunyxoZ9jX49mTM7yWBkH7qPgqNY7a82bfOiRr
pFKud9RUAhbzeA0FPxueY4SsHQ3ZRAp6DNJ7iqBJnTOo3BXhjA2e6XXVGQv3bUHI9mDz4uYxhnwo
U2MfegB6jZtkDiYinmlru3Q62q2G88GJiCVcGEBT7YOiYyIhp3qt2UebjREgoVE2ujJS7E/JMsUJ
OwynP1+f9BZEFZLd/CUBHAfuYSSGaf65/rELFQjFwNUjQY7an9MnPZUeXKPYMWbX+7HERheHAz4L
VEylD4tYrkAoSnNPygMqj5uditfWaNuxux23nOerdPnTem2BTFxcDUka/cy16Y2qmcXueFCaZMSp
tT1CAuxB1HaUdZ3Xuu/uxcqu8r2xHieG/r/XWYDnHPL7pxndYVapCusSOZIZPr+GlbNfPK8PTmjZ
OX7UlYtkWtqRxVQpM+mMsZm0bc6xlwg7JckFT3jsapWjSYoFun73lid1xW/lsdTHtanNQlmVxDfc
Ghh8FSpiZT+ndHBTFHLlGK/LhE2JtIievJs55kF5/IlA49KcYXAXxTrEFgBTN7FV7MYLErYP4Btc
kFKQIaSjtSCWCxBnNQeuUs17EiGvMndORmZfm7G6+CkkY5zDhG4HrhfuOylYf4+KFHiVphAMsAWX
+i9A9uyGldpGt2HUNDuX4rzgZGooGgXZoCgdfMlJ7iVH6HNYLGSgRDlhsS/2mWPIxrjOwh0pVRqX
6gjd1I4FmTZR0NncAg6chAOli5LZR95tpz+2tfIP4BtiUqYlq5nSHxJzQ0HNwO96d07dCDkD/Pnv
/HKJuholGgIUzKAwJO3eVAM9Vifyy2LykW13wCp9krFYI00yNm6wwYGRqllEp4XK8LeDA4N87+XZ
Vbcg2NwZa6UWulLr0oEI+etU0M/uZ1PVcWk0U/HCGnuDmFwmvoEGbvuNSPQHBwOu5+eKfacTuRmd
ixsrDR2mSwFn3VCiRN8I/RWfIvuqlH5spbSGEeNoeawr4Jiyks7xEGkz6is9nr8OmPlY1ESCPDHp
gZCcD1hP09Phy6so3zSKIqRjTCNPSDeKNpy7AuUy2G9j083xVQzrrIe5K0Jyzl1zlboqOvqOErgu
9OMRMSYQdp9tSt+0qUE6SYonFOPiHCxRfX9rTDPOczRopGUFZZUBAVPgcKepV3sRfH1h5ItE2bhv
zIBDw0C2TkX3DmaBQd2mSJRIoLU0SSIZ7WaZil1iMrezeMtvPdlSwizYxamTUPMqmjydIfA7oN7Y
Lr+3M9KW21bfd/gULPJY7D9hJaR7wcout+ACqAFs3VYbJnztOaW2eckSYj2E53VMUtaODAERycMN
1TblQQDBwhr8HNYqvoZP7vWYefr6rhopWZzJGM/lwEZdtl6T0H7rXIiFcC21kizHbcBgFrGuOXYy
ebX35vYxfxQ38+1xJhaDdaHE+iaIP6yeURVKSPqS2oslPXqxPxR4L/4a3dZ4iDrSz1QOrYI5xT3j
itboOHyvkzPTUX9iyFV5TOZKrjU2S2C6FNYWe6LPZnBV/K6pkMA0c1Yc0SAskPMOuHKOuKBI32HX
nnuNZ9jjO47l0LjrAdmoFD/YhcZlZaRfuRJIKKxPWg/mGfwcVJwuajr5SLi5YNtJ9WOkxr1BN1vq
NnYGqOiGZKPRIBvPru9B46L1qJ3w1hpgrIsIfFz9Lbee98PRfQAwV2yLp3sWeY4flofY+/WiFQxs
4sZoHY+1dGfZwUHKoPDaVoJnhaQMIGm9citQo//VkaZBMYKRixTLwQFbkIEc2wS2gzCmOec3Hd/1
FfB4g9KZ8Vpj6qC/0plUhWSNDuoDZlQbx0fjOvsRBwhqEjQP8Ym3N+XTPUMsv3g5NunFQ7VW+i74
ekhbuv2E4w1f+dkfyHU0HkSSoLzy/sS7rqewIChe98WTqRigSjA5EwMy42fHw4PM4tX7jjmtXoBC
IpFLqvqL9D4dP/GDhDDNf6gu4LTMOeOftPdUkeYo2npZsJ/FOjJ8pNbXSNUsKxF8HIi1FP7L76Up
of9U9DyaejEpM7FyN5Zpfgh3XJItbuU1U8QVLo5Bynu027LpqwOE1uboM2KTfy7T9QVYn9tTqQ4h
IVcrzZWCc/eW2mSJ8+XMysHGjza9F90Dv/f7QEV5bJqj5pFW/R8PbrIb8bwdV9A9fwX1vG72hwYV
JILvuJH2WVqsGikMnlMWjJwPsfUemwBEPCN93n6I3yBYY96lKvOR5ke2A1PfQQDl78WJi1Prmzad
mW/YTz+olBvN462iLl3y7/iIuoOkrUg/z/jbgLPcCOk8tCP4ACtcjuqNvthuYW2pYQCwi/Gzg27v
v2uEmIBkxIIfqg5g7gNZfcLJNSjtGt8kgGRwDQtOAerF0HUKxHnJf6BmlU3pjfvcn02ZttXznrB3
65WKZZgBC98CSe7xBYkCkNd33S9B6yI1PNWEI1SqQTc9NnDlynOTAM38eeOx8JkGqZqNK8TtD9fg
AlK6u8sekKPkEsbNic0GsVkEummdNa2sjVoJ84YDaY6utVr16drYFgGFsTZqQybpyHIJbpZs8mxA
Pk6blkq/f+66oX3qdPduV9GmnljbjMzKiLRtFX8QyPxjHieES5WH4WHSiwDSEzPZslIR/OLncIsG
A40dV/g6JDlvoaSLvRmoSDJSvrX6U4zcCTJM4pNDFhjLujEEMk7M35luHtg6Z57K1/dr24bRIDmM
HRUoNuVqpZrjVmSdfiB+3/0NC4vEa7HnyM8eouavw+DXV0eMTOd37Qw3I99XvoLjZVI8O7t4Q1Ie
JnzBx7naR84EqMxAbzjZeARpywkeiSm0QxK/fHJ2AgnRkp3FiQt7Zi9rxSt3AgA8aqnCmq713wsT
y9amVlxTiAP3NliBYNnpz2qhtKXh9kfs5uM+0gvV7O7hld6CYBFwn8DZtdbRdSLFZIueFQrhnrDq
HSZXkrOlW6HMyzr4sREv6L55Y5mAwJZFYiEV4xD67s3x/L2YqObTSkV07cMoZcD+GMfNAIdj3zkW
pZ84PEQSKzC7qomcoA4znAJkYYFpU8I1zMTDwR1o7a1eN7ra38Rm0/KpnrDpU0OftlidQ/sb6w1j
It2CWPkKwa0Pi+l9FAMovUGxzokdOYlDG1C86rzgccnBcfoPgmlrOC9f8koIGWZbYThHLQBU7eUX
3xyZJ0YjsjHYM+r6n3PLgsiDHGmmx40mdUbG8+Sa36q5P+xjMngObn61GkaZPYiyUvalexQ2U2hf
2nZqruGlJxyEI2Qj/dpvR/WgvlJSZDgPxyL/OT6l7gmBP8VYdcRPoomFNeaW1xd0ITP7LUuiiOEb
Rwu0rnPrEEzN7ZcPibA1ginlkEw0qTTyl89yHGodHo/N61ll2X8ls+rChmkPt15RJrBCAY92GKUS
lDD8hTwGDJvuZ7ahjNZTG7N4YCxpaLwNu0XO2zcKOAz118rfyGvLV4lsVJzQlonLS60EzZ38yT1Y
T1xIBuk2YUDK4CjQHFCbnm34TV/Dc3XyQ4fIn0rVw8quHEOWznTKREYc3VcnCrHDY2E4dUat1LxQ
gjDIobOPVZD7cGopjLAxZbeymeXfovvbNlH0JFvIrEQ9jVIbw64hDxEHHD5SfSaB7plwjTigm1kP
TtUty4CiRhOslZG3A6tRay5r4i/3PmfV2rHTTj90keYL5pEk/JuoN9gK7HkBAlTluBhabj7Qqe9w
Xs6/8Qlmn6ZioRXPQMVF9XTetP3lU2Bsy0JcpUzwuhiV3fed8SPDYoxe+Rux+m/FZEIj3xERYfs6
FVa4XnyDhgynzwjER6acRMse3di1oafMWZUF9aA9xMRMzaEXM0goZLPYjLXQMLGOnH5KuQbxA6mx
xJdm5mZX48aDKGEKIMwjjD89Us/OB4cvMkrgEjwBNZWFvNYoca+5bYeNMzrGc4iR5JyVO2rKJhFU
wG/xb5xEtIUkHMhyQNM0l7A5JbnxgxNeUqGew8Kna4mcyXlcGn1lk5EETZHyWW9Yv+/A32UwNzen
kMaHoI1ThUDLDO9NO5mIciE/ADAZbSChEqQIad7QoSPE8BvtvSKhZ4uPmxXo3L3asgeMDKf0jpgI
P2Bxj4s7W2Wo4whbE/7Uhf3e+/n0cxkZcnpJwhaPElw/12IBjWenDl6udd+iIt4Oo+rMMGK4z25t
GL2MNy4vdhHRgnwf9Qw35hL8MVvvnTWFiXLNyHO23n5jWBCHLucwnftQLnIfMb59B61+lfycWeKs
CN3fw9qFKun9xLcq/YekcFeAK/i79ddUTTzkwflNjZX5rktBm/WdfxWKyXNHtib498y+vkTcqxCF
jBgESS4shTWmRUZguHKKnGLy4ZGS/j5evH6brCtbc76d1RlWeyJkmH6UnwngTOMvausKPFJfHZ3D
wa+ilIU6gfIslgEmHtx574HvL6PwmC9y3H3mp7zefc3Rk+3tkro/hQnQ2o0uL2RyxXAA/VqhWzOL
1MIGauHxxJWedj8W0SOttqoRd3maI/no/nMt557xV7log9A/JO13IZMR2IL1br9otvfRSrf3wjuk
1mMGClRja8jBIp257T8ISwn2AND6nhgWZj8sRyCmaWO7ot9r7wloaeUcJzmORHC+V3biexB9mfkt
4rorq10NoaU1koJcus7SxQtNS/Mf8rDMn7e7MHPOnl8k+ktAAZBaxmquLAdjKkNjTcXaj1cRhXAi
oeAgXTqxtspL9qZ1tVVktRLWmNPtlH9Do7mEPy+IMQDL3RkIQLa6705bUxKq3BKYzfMManXuR8GG
3JFWSprWABE37F17PgqhD2rSvtZNNOnFx8Fyhj8FQS7j6qN8oNkbKy8Gsjl50nl88iYzS5CGul1t
vwXrcGeCiS1k+9ek3YcXG5vuN07Cck/e+quo7CPu0btrHALzCekUCFmAooRSiiAnMbkEExiO70Ru
m8GK2RhBpcZnzmV28t55jiCT5ErsCxMlSU9gcyaH9MFbEMyiTGZTZQUlO3eY/i6RqtQrXZnvrabM
kmC0zrJzVT+Utc6LDbCq9K13v8XwI1PvAVbn/CmVx7AkYNPTbUGgGNrJIRNM0QP5HbEzi/xPOSF0
6WTQ8lSCctl4n9gSvGVq5lG8jmRwG2fS8dFTgSj5qMV7gmIWbZ94RGtRP0LBbI2WPxdy2B2MAo0E
YTgN+D5ZiBSC0RjqgRpVyrw+E2/vCYXkockB7RFpLdeTNGhIKP7rkqEHIXnmOpU4Ob0HOwqJUY45
ndacAi5mxtm8YutKcY2ceX3+MgY8AYm9qnibhLJQ7Z8x92yqXwEgWDv5niNSRckEPyokC9trMi4m
hDP+hD0H13u2X1zD6zk7ZmdHtIpjk3gY67N8w4LjeBUlzlwdHPe4jJIX+d7QoH3kab1dSNjE+wZG
V66Yo7Vvz4mpQeOi+vYPcUwozZ0cwLwQoDwKt4l6qe17yDp5G6HhtDaCSIPXbmb4Jww7GYQ9OCdY
R6XulAdv+u5Y+z1LQ5zkg4Yk4vdepXq+YdJ2Kh03cOukXAQbfGROS/Mw8k4QH5UMLo3e4syuEVf1
iUioFqzohJeJLK8wIaOhEYAWZNyXKpVGTHnJQTKVnK64L/F1QoP54gwc+0cpBJAeyrEPQn2XmkT3
GjvGyOaoTE7JybRAybYmqdvCmW/4lb6uaDwXHCx4shp3A7gkZDSbOzlvLODOAxmWKqAth+bITQBH
BsxcySvoO3likbKCD/XFP/q5tRcEjgH1FHxrXetsx+LSS4W0PznEN83Uii8EvUpB8Ewz8GRNtZHx
mT4uCw7fiN4YvM0ftA1bGQMLkq0B7SWABS1wz9edfTJzV+m4K9FxcyyAyVxSmx93SsxPfzkZHd0I
5Ci//ct2nr37xx62CUyk47Xo+z+z+FDe6YTg9XSC7OP7XIYHfyt+dPkzqBFtkena6k5FMXhs/2wX
wIjYDFuO/HNazMJvQAa6GP6e32E+tm9ZFqYJzR1hn113NhbZHNV5ihR56Yh0w9tBf5JlrQGtpoq8
Ni4GegVzP6ggcjZ+z5aKGBSMm7aXfDkz0aYmGo23UUYrNjabSD2lHTCj4KFGLQO4FJo3RqaTQuyj
1LFY+ciadeh4FnlMLIquWJe1gxm7XenHqM8Z/JQT9WR7BlAN7ct5tYLk+SWfHYWyGqHI2/+2UZu6
UQ3CwZJlpM7HtkjYvADUr5cbeJ94Og4v4Su2PMR/ST8QTUvwn5P7NYoE+fTEPrisgSaEpQyUts9v
wJuygavG+9XxaNtIetJuYlnAI0yeqzYsxks9sjgsxXmvCvSE5d0X5d0NgLqeIoSzpqIs8HNiia18
TUgZB6Lg7UyUgDPf9Fyag63ZfAuyOE2vmkhtkwnTt+KRRN2/UeFm2J3/ieodXdcBlYMxOKXoYnbh
TkUetRHJqlrp8aW8TRLfLo0BhEdyt5ChU/FMQoViRBQMYDv0qMEtjCzRQUcTT/Weqr2CZB/vOby7
rEi5qVGWn0+Q5pm2+T/HiBvDlVc7zamQyYQevGMToTN09eK10KLVwWXd6snFE8zwQ/ohxS2QXlqg
n6imx3m6YTRHFUzhXg7Geisd4rEibIRAr7XhaS+oOmaS4DRqS4ODdJegaZDWXrsXn53bJeaUCmJX
ILw8Q6iDAyVVDoOZWkTbC0WOYX4nM8G7C5YRtouV6TSwrhKWcilaE9LLjWH6DmAuFd5A6YZaiJKW
yK0RxZM/+roAabXIyUeUa+KnJXxXQvueq0Gs6cZiwJjMVutL4VhsAQMZhducCPQtQMXfZXOdlBfC
XMOp2+OZIOITUAdeF6se0jo1AIsbd6BxD27eo+TVkspJiwwmFGd/jr8PUUvh8U+8YLFg30Z9/9hw
0dncn8bt6M/P2jGkv3M9kHQR/FvGIEleqyTZ3AKm1Nox6ieeQg02gK8Rsq4Qoa5uopPomKidyd/y
DnTbGhDhb2+KBWPryQBTM2MJIi3oFW1XxmW2ijcUrlRBmJp4ufRUzzs9pCw3GBHYR+kN5eZBqVKY
twR6JIbK+hH4x2gwVYr833PkPG16YlkvaSkDfB4TYgpzYg7MbdXCSHK/cjem4k55hA/66EX7Yfin
a251MBvHT3PmV3IHJ6CbRe9TguprEafSd2fOCf9wyivVZ1VuliLEtWVTDycwh+/XAZGWuTpJBxR2
UQ2EWDkbEHeJANI9iBwMgyVjfIZ14MMM8lrlSm0HMYF+hpInYruFj1tg+5mUBXBYuIw+wbnxCg47
AIp0sEEhQD1Q2euitRixitTa9+ToyuHTLVBblAzI/5iZsmX8Wsc5L5WLYzWmFritBfloOVBUYkmb
Ppv3r7rJi5pR1Db6V/b+0JAgVtH/CcjkQujmBfPyKly/dm76YRTK0NgQS78lHARmwd0KzbUaiB2J
owkqeIhWm1PLC2cHHn9WYbjCwh/qKkIa6as/q9tLTyOe4yQO1UE6woiDxQL+hiNK5AV5cYtgqdho
3mWFKSAeW1IVCuCp7AvzrZVN79a/mF/JsYUiYK9uo0l17KW5CCvO1Ipgb1a9Y+XfEhoozbNl5RKL
Fwm4TtdVRDSQ37tC4CdK8jJwNdpb0LKQX25ih1uclsvaRFaivOEedthboPJeEsbvBb/9ySmvh1h0
+TjLYrB9iGdpNcVFOMYyqTUvAG0cz/6m1/BA8ogUws81nACPmpt0H0gYGzaQJtY0ur51nGb0nVKE
Jp3e7p6Gvp20JMfi7RlbtuEXuVUw6fii32YwuyA/1kaPKkjLdG76bgBkr+cHID3/RwpRdGVnwh85
Jey7Yt5sYOQ2736/YbjXRGb9gGntWCrk/6jPL7/RMiYrfmNStBRBOCl1Tn04vwbHB1kko2vemeHq
tSz8NkKjg4IycRY++0waH7EzydaLKrR+TcNoAbPhgfTOLB4cAxZhXnGJJvWwAO+Oup55CmcsTj93
2DdUcyT3nDVjwuMhv9LlY9valgv0SyKYo/ilWU66Vq0riuawzuGyKTixkp+2Y86u19TFMsgSJg1f
9H9bnezJQWAOiK/OECH/qWkrkz3NwX6/Vj4dQ7PtdM1SbR+ybH8RNDfLZem4j/dl2CYtPXzVkJyE
Qqq+rssoL5E21+T3lm6JL2OmyHrjyJh6pv3MF2bY00GjUB9FMWy2vDtR9Niw70x8wImPAuKYbUtG
SEaYzaPrBeJkPe5Qx1u6RsFLr6NzIUllXGJo4a9T+bt8FEOKr+50kQ+b0tCFiLzCdaZq5bAfEekh
IXP4YN7o+qUUmvQG9rwuPf2o/hFnKHk112WqiDGtvBeG/Y2r1CL11j/6fP7pmltPRYF2K+HcCoKO
IkG0MveEesKvjdM6N4PnUZe6KcLZxRwTJc0xTZ/L3LYXtwCD2OV4w84a+FZGCPdlliuRrH+O7W9H
t9Q/RRwyh3ObIZnrfMsLU1BQYw2HmzWzYNuKiyfupqte/Ood2gbL3xOnrvw9y7ES/UdHn3eo446Z
zBNi2pffHSZGl3/J5WAshC8XdtTnkYjG/0UnvQ/+SFMCMuvIWagYmtyn3WU3jZxrN9iqwSPo8h9/
ZcFqfNIocDjYNWTojlUm7PK8hGtatAUemqCnQTRrhqAiBq6ZB3JR73rYbazK8B1QON68tC8K0BxL
g7EDPsOCyvvYlm4Zf9yBj0vt8YMHbL9q7JV/wZcLZhmVj+uqsgsjQHld4wFfvAcMZ7JVpsaerES4
gQlznZ/XBWZrswVfKXMyJouBPQrDX2/6psEL5Ihnkr3nXko73gs3YEk8IxDoqX+oAMbEnLNwmZ40
CBN26uLak7weMYCw5h0clhVcgnoewiwdhkL3cNgO2SlUu6MgSyQqLVzpAgXIoVQpqZ6CFZyEQX+a
XubAPPhdUv+iN1l2KM0H3DgBVN2beWxoGwItutJUnZL0zK2p8Y4sizAAXDCccc0axa6hA5GsBkFS
GMsHggw6kCqI+6FkBln45fDY+3RrShmeT5ess6O7nUnihJWhj4OfGv2lCxr5bx1CW/B1nC5Qrmyq
E8b/wf3K2zHOp2XIP/NGytlxhx0JsQz8HRjPzr5X2Nv+sZYJRPSTbe+RX2Nkjld85hT4ShQzr3z/
gXgAOpO7w2QoEdq3f5xkLXjR4S+WVdO5NTxWA4H2ovtK3a94tsYHxffSP6sBrB5JayXv8r4Taf5k
JJuS117SDBTj6qjm3crDLpmJVK4Y6YGqQ8uC0um5PaukS4966rJaH8s+Zwx2PSJK83DXRMTCsEBl
W9V3PfXdg9dfJRuJkXZDrZGFNQfXYPFMSFLHEKgYzhgXQVUXdly9oMoqQrr0l5EuOQlzRbQ3qDCf
vNKKm0o73gEDlM8SsXDVWxhwaUiHjpzT1FUo711gwwuy0JbOaGZYwXdUyNbPGD2uYyT6ijbMkqgw
P/nBl5YF1Eb11KJzowv3sIKUJJ0mGkSqxcbxNLBvjzdyfYVzO5vnngOKiYl609qh/TfqL893q238
iYFovd5TW3EXD0W+agXfYHEmauI6xBR4MDcb+zM07ToaHlinZoQh3+1+4EJHaGXQNx1ryh0c5o4o
qxxV8Jt3V0HsMaa0W+UgyrFAGLQ3pHkT2MI3f4IgTdA1ptUReIiApoH3n/bsajCFVljZEFfPAKxp
BoUg2c7phngMs2lFZ0tRmi2QYvHSNxeQ2UOnAC0CEVL4SDYnT7XY6Vtip01sHu+rXMISOPNUPKyE
sjX5PPsPxvN3JUVIT/wB95+QSiu5IwErn6Wf74pqVuv1ZLtgwevROXYX+ytK5Kn7yOVQ8PiqR5pr
GJv+vmocxDECOcpTLFV5+V7LcaX2A8EggyA0QZMxvw98LQW2/sC+WgFioK1nX+BwLrlBkmbtnJ6X
4eZWA+m8eq8mMAq5d6xbUBU0bov77Mw6ferUFVx4CD06JJa0oCTZJfA6V4oDEVCZaRK7lpK8Y1Zw
lCIX1Vnns8YTPX/2W1IryPSL9Tua+gKLWB2DO0PSRtPG2KNccRY773MwOuMDUPClmlIHT6yDtvuS
vZxjty8f03dM9JKegy1QJoIfg/M+WQdUbER2F4VzrpD4hpCLniocEtmPSBZP0HyHl4J9Jp0iKSLQ
kWJjyf+lJk3JA612EcFTxD+mJtmHVZeqZhkQUpe+LL6hsuaoFXijXJeobKaJKNT8ONqXPtnuVnod
VMVh5OV//5FMHdFvGrI7KT8Rm6hR+198MILVXvymFF0RtG/ndCSl/Ta6CnQFi4Y6Q72OQHH2ZHq0
eJ7vmpaMNrWByyXM28k3o5mVWfnREny6UkBxbe7fiEjKnsfRT8V8c8tuUhCXACC88aegEmsCYmVs
5wXoH8XMP7MfDKWumVSNALSnInZ79WKXP1rjmmzCIUPkU3agyo5AUsytJxc2SwF4f3fip24FeHEZ
cPFk90MjWj4u2uBtEht/YJiFM8MDNCLgK4L1h3VGko/0fSFgxyIlti0aTGWVEK7kZ38LMmda0aTc
7F53B4o08SWvz/SnGgjIzgxp/seSAkBhPiqWV+rcfsosJvll25DqLZx7W8F1m95j3Kuo3NuAyxVC
R70u+LOMH3aQ213/u+Y/3+OZaGvqzoi7sZIN+iVzOKtdWz/Q2qsFEkwQ26pCUs+9GDbcotbtFKaB
JJVEK68zPXzRL8EsqDK2DJSyxrJUixEgYx0DnSOjwP9Jx5FPAVewc3prk3U30AHbAhzVCdmypUuW
HSwlqWyVzces253CKleKKDmdK11fFqyM6ZD/LCBJ/iK6N66m6ymlDCDwsbfLPM5GyRW9LMk0Z0+R
sJ1u+7ovDYR2SVlDz5Z77BGMEUJXvKJZxhyJjbkmYsWzgHOUDfg1b0XRN/bjr4rcO8KX/fh/2Zhc
a1QMCP+PI7xpMfNFiBnh1TqKb2nna/uuFfHujG9VfTU3Uci/Wbc1h+je9nHwsQ84u/0j6zNwLiLo
/kVoBJQFS2TdZUgpoMUKKIvalmcLJFDzs15T6pbGPdzDcUewPxR8zn0Rc40zhXFYFn8UuXuaHMWc
kON4tPrhYIvWxzRptq0dvHMRutNbari7sDI+xUpEsbKMRVIXK1IVU2ADWbIjp9BsNOo/gZ7cV0rs
PVsG8YgfvpXC00MQbfBjufpC2Reem8A7SG1UkT5RHnKhp3sVVZmpSpYrM0OwozPpkZ3cvGhc229S
tgyP5na8JMABRelIoMwq/YCF72+Hq3x2jI9s8STxAIEYripmqFKRSkk8yCxrGzDAMRisBjSVro9T
7JvQ11oIYxgYPJxsdu6kMCcfPEnzlswIJaC4Fwa3VGH3xUNtaaADAIpTmZof5/cGtLVjCjp+Jid5
VYvWFI15uXn726kBKLjBInYfgeUz5UXRnHpDbXrNVcM2dNtbjg1cLajzenJilueuFfc5umxUtH1D
AJ7V37hUV+CV12iq9uGJd1IqoO7Cde9MFHrHW6F+/N6czSrf7JxrzIK9FOzyS04I2Dd3uau84ixd
odYAW6klkzevZG+x7EoRs8GR3WpdyBx4o66hiZRQmKHajvjdh6ZJFaKmuHweTkX+a5C0blewqVVk
6QO0A6VCFI9Px3l9l6XSZJZWpIWbOarbMTq5u+vAuBhLpFRtuKz07YVuEGDcIgzUO7fNRxye4GHh
lz7/6fklA/BBRAbBTOV2lOvCFdd6Bm6TUBUILZxnFOvq1lIDhy9He6sMy6lFvOe1tyx3VjHHDGql
Vo6LSO4ahuhhrlur26E8WknIbejF4kz0pQgOUvo1/HscH7c1KycCdpGuZJW7Ktywl8pTglXYmO0H
d8WVUm0kHKFesvSar2y5/Q6SH5hAML0vRYTkttG9ARK0pxLpyp9+9aN6Ph1qZrisNgfgfZKI3t6w
1+/BHsUuV0FnWXmH6Nf/ByWIILObvi5+nGnoGNrmCyGt7QXK0eN3y2lXlG+qQHDc2Qn9H3tf8RhW
nXxpNil/Y26rPm8QkmbXexG2dN6/8ktQRI1LfN87lG37caZ0WWlmzeAUySvugfdRboVb1BvOcYpU
q4TNiuoPBftcturgHXpPjmDYZhGEjpH8jHjcSIlcJYMkrpqTZxOI05OOvsD+ciCWo4TxlrsTrhUs
ZsjCDvTjDa3dEMg/p2tgQUlyTCwbW+y1tFOZjLDZ3bPKyRoT0aqo59U+xPmMSmMZXw6f1D/LWvRG
C/EbNdivtE6K/SMP0dkfGYqDILrN+KYEUPFNVh/8EpMNUPbc/wtuWvEmW176KVG0lPZOZ1xtc0Kg
Bur3MiBEE4rfvfi0DCjZylApBD8phqbDF+MAlYS6wJgjrsuCEw9T6un4uFRzwpYeUP19HJgQPHGX
3D0llyK3DjTPcCobSB/Kp1XDd5MN08N56WGFzLq0jfiXTQae+xUzvsmYQ12+m028Ptb0o1+oxsFT
EdHe+WmgsTq9LiqmNyW1kc4mHHCF79PNotrP1meiJZsM6wnHA0WTymrCiTcsHqRYKqFhlXT3J0Vi
r+9v/yjWJ+DUprIMXdDiNHBAqIY40xkewljZqrHyhp2o19d3IscJmqyDCeF2PwahEFweujWjnX+X
1p8SE6xAMpZ7BPQmcLe0AEnbmRJWjRx6XQ6+Tkow065s6bk0HMTCeDyueIAgAMtBhTu3PquNpIPK
pB5UIM8sTg6V7gUYiWe5UGMVC/gNA7H79XFlu1Dbh9FYS+FB6PauKhAat+/odFKbQREEOv5x9/jy
QWUIbGXt3gsEthgg37e9GPyfu9KztTqa525o6pKvrkLnFqN5fL6F7Fv+rQXqRslxSHfsR/PexXYF
t+rZfU0UeBrEWehMn5LF5mtWHwndW5SZT7F7+rmEqyMT/k4c68mH5XBdZmVchuQgGpxnoaJHosUn
Cw+11Jkdmz96Romur8WPbUhCxRZ3nFyvNIP/aoyc6OEBsW6Wn5csK8qnsPZhMVFeGpt1yHqd+g1w
I2hpO0bWHKnXI6eQnX2SRqgWctbbqnukU778c8XplR8UEVwzs/LyicO8l550z0OBuul2aT7UE1s6
WhC7upobZHNvJtF37tpfAAVrSAJ2dire5aVwV3lxTUlRrOqFv5PQIxao2nfm7q7CoN8HUyXtgq6Z
yQn9cEjanFVE6b67jN587ykWSWXnR1PoNwx7406RYI+DQtajhXV7uX3DpDXANiNTau2mkwYog0UN
2hqTvdZc+Co/V2ylL3tGZkBZ4hKwO/TU3WbkD/t9uufhxxuSoGK/xebZmCrXKIBf5CXaXzmjyTYm
zvTk6fvwDIgGKw/KwTPDsZMlZfjAxQ00a2ZWfFFgu6crAEQS63cb+YMovDjcoENPLxw2iBgGvW/e
Kuui9lJkU+8QuxZJmqnQuUOCNZfgGLIq7ef+Yt+L9hzXqXXwhfRboDmgdTS6zA6f4rljg7OOPo1M
ULaOou/xJAIbP16mDm21PNVx9yCpT7W8dGXQZgL4dQ8L2QQyV6lokLs66MGr+dnRnWxq7ryCRHWW
9mtGIvAypIW66bjhKLdinuPANaAn+noFKCLU1zd9TuTuYRQikxGU0S7paUgSuBnyaQoaKkcqPdo0
7YT/A5UHH2He71chhSSaR6gumVzNIuV7NJs3wbQ8OK4uiIl8kMliXFPrtAQ/e5bPHDtIJra/Wlcg
vsBvLHA5E1xcbJ4o63jffPwcJ2ujcYFADUJCC+M90YNWk3jC7n0qwDo29UIqsljq2XgwRpJSpTYj
KVsEIngFPCvfKRp5PZl8C52PnAGBuvaVdOk3qVWY/4nN0eXqH7eJTAijFj0zUPL4mhXq2TaoMw5C
f2D+2E3DS6eiVepN3vxp0vXqg68acWFa5U7cyWtIe37k8phF8bXNP+63qH3l2EJS3dawHZ/GYx9m
gE7XWGDnwcB8EzZt5Z/3GU0MlfikJEf1SkQXaWQU4WqMln95O87+hHGsWzXFdqZCMlcDoOYJiqiG
er1rwrFjP4na1k6sLlrXFfVMGOuWIXj0rYE5XFnvCtp9WGAW/5PStQ1+rG7kgF3pS4nCt3ne/oD6
Odvf60czy/AGTYOPZymLMwhPvMQ5oiuy479qKIg2T9/bHwm1BpcaP+Sa/EipJeStqtqZFsKV3YbX
7ReIMfpqGJj6yoCIcJg37n+4kWqtctRkx2+vttcy3kjvnSmlpkZbWVJTj+3xpwpWALdpjBPsqT1I
WO6BFIRgAZdSpiOfMXpcclPhtCgxktbBESzOE+PXQZ5WZrSHcZVzLIDZZbEWdQpSMAnNW6RJL9vm
k0EDg6a6E84bMIIk4S5Ra+YEGULAKud7N8uuRbG55T78bKwa/OiLr3vkVrdpwYywounzxMHudlqR
tcXh8VZa99+CYSpqW8t0VRgo9GfJI+y0gDIYcdOooK5uCZPrw/9lGb4v1gEhVadoLE9w7Kim+8lE
uOzR/nz335Hz4uS4FBlNsiX/BXB+vwKfBCuQNxLjnGwPrzKpZyylVggljE/H5m0PesZ9ZmCQqrz7
o2hzMtzwos+JhJUk8O/ZLvx64KANpKBRFQUPKfy8VWCe6eqfqMKG7RbsNyIasv7B6rE0t8gSekV/
7seKy89QlhUxyjubEC+ZeHc0RMhzdmvrzoWK2qdS+xmTKUrtgKrPG9inesw0OF7a20ixSm9ECE3l
AjGXTzFyHRIbfKdWj+mFz/GSNWCtkzUNybai8PfhdOpSSur6repznRpiN4IkieSKkqzpK1bmyPXH
EUkp1jsH0T1xMG8dETDPkS/VFmUkbOiA4CMtrNFdMfemyq10m6bPwCPdbsknHoelgZ/dMo0bdY+v
XckpSmozBAqiqlST4GJcrPwXSikoFNl/li5s95WPqWbOl8N8sNtY6IOshWPgBvRFHHpYeTZHIX8m
HmxycRA5lgeSZWX5HlOhFtudHQH6NlzCVXsysILnLUz2l7B4a8CZjHav1Z+KoBxcmpxj7tEypUtf
g8cVPUEB7ZsumSOcqrfv9UjKEvFDWeIiER3ENahDJnZ9wSwFXlJlydVU4LhT0hoHG1pjoKfKTcnj
ItWEcK+AwdHf6l4RIoz2MS9K+M2CPDnBkxrThl6DN9OVujMTGIH7LmhMM+e/K+VVsfZPTuRdZ3ZF
dXmvdCgDORk2ZmNAu7sFczboTBPhJJ21UOajuoHwe6mIbiftxzXfxkhx++vKyeRSCp5HdoYlimbm
AAxKfi0nEdGr8mugeZcmR4YxvVM4k88jqh61cfiWac5LzHUaej1JZl4S0hyakpwajT762lpSmGzs
hAPO+WWoB5nJEkeVc6NjfCcNAEVH2Kzi6gxLtKyt438MD2iSFmgXjiarxNrOlFR2NohbiVxmZ/Lw
GIFmkZM/ZJIoEDNtW1Zb/O+CgQCezVX45EgqPiJAZOnGPzAdZoEYoEmLPC1wZjUU9dLqUzR4qS8I
3VITu7Rbp9AOeKC96OPUpeKFDnIDfUza+nHVN2kyKEKEaeLKrgoKBwLUBD6hZ6vACF839D5RqyTa
MFtGjtvLlkH3Mjx4TT/092g2THSNMiD95cvR3BJI362xEdfF4LAry7eMGog5kcp8DPF6mvdwF86p
PDhdJbUYerJDwQPLm58dNlXNdwIiU6+PrcKVLJxtzCHADVwWxxGgVkKMxS2CX26H/Cn4RTFOD0SD
73R0NCuZoHY7C54hPE1eAjUdhyM4CQVQw6MvoGI8fJXqgYvCdOTSclwrB8+rNLAEHWuIChW5AS+V
nWqN+KU7YanCPWjEQwk2VNwKdl50uHjqKpFUsikgtWYESDO7gnkul7nqGxre4VIpweeQEydVomAN
hx5ta9gauEUwudHqq/8aMRWXJVtajPLDN+vWX2wPTT2VbfmhUYrOklYAuc+NUFWh4P4cIqJHVgVG
5f01vcIHFJJGgW2F5PQzFD0p7RLv8Pfm3/sqlx/YHvotHW2c9fkXpJq+lzCQ3iszKjc3AVXSrCGe
63JyYK+3Pz9fr0CQy4x5qPWrcEGvFItLGx2d+yilzEublkT0n3c+I5UrylMrfC6x4AAEPszxA9qz
FqZJ/50QMV91p6eDPLjExL3N9VxGtd4BCqON4hh3i4U49ftu0P0aiCv96x6C4a358mIOC4DZhtOo
2+TiUiABk/vGpFORKJx0ffc1S/WxIj43SjeSikXuszJwxC7ohoPQOD1VkHRERvHJIiBXA9293jou
qDTui8gMYec5FlHN5kv2pPIdnW+EaoQp/hH5EY7wqXt8NCf5AVcH0GmdLToT3u4QXgaN42j+Azqs
XNvvQEIhkhZYPK/OixBnKlXmsk+HN4+7ebNiEk3Ad5mwztneC8CXyiJqNqjI1/B8Un5Wezo0zidE
wSGtbxuMGvcfxWipY+j03KmN+G8UXuhdShvhApjxD/akwfsN4Ak53s5Syfwqh6m+rNjmBSSie+2Z
hZRX+zcCgiZz6J0rY8XQ6AHum39c5gzzbYTvHt1rZCI7oFh1e+5JgAy1Z8Khfix2U1utEaOq3HLr
WrktKiEMNEY0Y6/KamWZV5whWWDt/qDOUD1q4V0ycKbyeK9oUaAXee/RMivzoXB5fYlB8ogQcr02
dCXYPyvX7Bxd7if0WRZwGm7Xyi35SYaxxAyqqcm9j8FS0vJerJ6AAX3BTMWJypSHrb+9bDOKp4Ie
LfiiB6mH0oGzCe7AaVTLg+riKqr0VF+uWljuFHcdBy0pcy1dQYz6L2ZCpiRZwvV7RC3zj69F4nap
/bsn9gKoUexDz8xJKdVFxYzdcl5cgxyTp+8zlmcAmvkDdbI4PMYH1aNA4+mUZ1xy8ZJFOuDfyQO5
KB4z+7MYrJtbQfMl963YTnkaJcd4gmbi8dTC0JMm2TSnA28TOLBuz+aXoJsmLDOK28fSK8OQeWyR
S9gci7T4/gapLnlb/fAJHlTNLibhCV5VTA/bykGuMWn5DDgU+vRk8UmAFutQeoO0WGBgXM64S0bA
LtNGoRzIj0GbFEEQLrmm6jqCBK/tCIsk6zEaRfVw2VBsJsinQUi86N4JWMcfWFGsSHMgeDDsgvl1
hvsqBc4eQBF/dqcwY4nT7D4HeZYltDNov+cK4nVyrLU+1NQJGoY/G5qE4+MgPD+Ml/ScgIU1ovaZ
vsb7sLgjASMLMKE5HlnqnYbUT0s7LfVMxRITlHtSgxAwJdHwVoIsg24qNlHElMgTBr1enI+ata+N
FRnwxeJIQguEPdxm7VkpaSr4JdvnYKSp9HTMB9tNlpXEMQbG9X5eSDShzK39qW4+km05n+eKZMZd
e1RIzZ7BpD8SJV+mSFVcJj7KeTWmKN9WS+TapGxkYh20BvMFMNLQ0bFl+5aNlhWEFbR5xwvtIM88
7GHloD8y7g2W81KOJdXuQ3WU+DJa4aJcGPZ8yTusQfNnP2BEpKYkbFV1g+N0kDOjlidb8WwrJ95F
In8g3Xg4fOLuiMPZ/1PYHFPJD3fD74YlNMNGo3pbutm5Npu3Cuzw+SfOz5LFBEZHOsrzJ7EbqljY
L9YfPqgs7SQCv80xMgyIxVPiS/kb+gP8WSFtK+vkdXAP9T5RV8P6KLFQ0/e7zClGlejdLP51N07n
p/ZgRTyHKiVpSL+GWcA+33N5Awg5K1OXLxHAZf+0fDDgrw/yF6n0W2G+L9PDRkWohtLagFcwCSeb
SDjPd8x99mkQW4KuPuZnKszuH2KC0FK3XdlmZm3CDQIlOVS8/eH75Q4Bp9tmcTiCLqJPl1kPoTHX
FqP/AQZpTetB0Ol8Mg+FLbt0ETXsaq/0F+0czA9dO9P/0zvulfi3QlKFkXD4NOsqxrfsrnqtcgD5
wPIb2iiesGk7DqnSdgfLaUp5JTReFnm31fOVS+cUzgkTCmKzHniIkEUctWSlLTqFHlrzev56jP9v
nytIC4qGpU6DcA6U86caPj6ZN7JgPgaybmKbdhgHSNHfhVBPevC72/AyqYcfD7/wS79lS5gOopQj
vbYcupO3f3j+764/zPik5omrPSkoDXr/Z72KOpAuSZexInTqealE0PwfotKrB6yNAP8dzA28m+vE
mwXesOi/WlbuC5GHxsbkK4Uo51qUyFfut5fjE0Vv1MnzHYcyOxouXjiPt/KvQFPqOZpAvmuWtkrj
hlYXwNG2+b/JXAbz5flsF1gzBSJFNakZosy+LITuSjGipq/lEzG08FWdLbVIXZD+zVfBpaiTlT7Z
D/Gs4XKDqbaeofUcTQQcx9JLM3sDyTpyB7zL6XLcr0IxmDhF37zFN51wgodf2mO1neuvolog/qh/
1W2SqnZl9ewyRV9UQ2+H5B8pDGXuw7pmZuMgfT0FgQbbHkhB8qvGilAX/o7yucJl3zDRhUGfF0c5
rPYm8kX+/X7tOB9lW81OWxHdxB2wkLBOzH3L+Fq7CHUnYT0eR99RSgmnHLunrA8ofqswhy4ihW2q
KGcsbw4y3fQojcQRoQe9qt7iPJSNPTP0436aC5y1eDEkeR2H1emX/Z4sy+B9PEN4OuV71jm2qci3
U3zH0D6C+A+nfsXcMqainznLDiQGuWR1RNjwTRRWnFO8D86gSx2Mgwlbi1//7dwd3t3tWPitD3wt
VfooEYAYafDdluQ/mPaydsEgpn9+t5eMOlo4FX0Jl1+6hl0/F7ExFmlu4Q/QwO2H/J9T1WnhODRC
wO+yfIPLaVVrI3vrrpd4xC9wiMDQ+xQ/FVmrybU3D8fx/rAVGYCjgH59vMezhA9ruFoVEYiNACbv
eDNC2E5qPW4jymBCIHV8sPnlo8wzp2G4GmAZdhVLrTvfh6WN6thpyjkh1uCmwUIPQtf6wzpgRGp7
zceS5vEsW8M3qRhPwG0gT88pwGRs0JpWT8Hd5ip1czKQtjNuf6AKe419wSePpI+rl9nzzdQUCe9+
tDUdRF7uN+s0xRYl2k0JOMVPyP0WmXs6HdmvNwtbFEl0u4KxbtM/9AHtpfKniHyp5Mmsx0sRU6vd
msPO9OpuGRmUkZBvg5vMwX2prOeb625ABchwb08ICgicNs3XyYNqHWkodYT8NmqSZT+zCxA53hla
huLtpD3H4Cw1cZeitTSOYBYrtVswWpK0ImuvtdEVUgIl+qME0NNgqe/wXuaHd8qPjoEk/QdmHnZH
Bbg7AFUzPvIXyIHmfVVGA/o4FrbmS1x/ZuBF5gsOU7YfqONAQaqNVhaBDifIdhb3XwSqNJSuZyLJ
C14nP2/bJTzblPoLUCHTfoLxgYWQZKFL4do1VZLdPtae1fXkDYFYaX+wW/dw36NbJPJ35IPAv7Ax
vCdfVR4y0k/gfyX580nvzkOlJ25aCDu2h1pFozHviNcay2bM9rXIqmUZIBFTgM4TUKnKODDhkHOc
AVzBEkRrKJfNFzK7duCygO8/c5B8ADqLvgs9YvEokTyKV2z6eDMbhTLLCjKD2omJsyRUZ5qcFc1J
vwjTmc8SY9v3uhJW5idi8e6vAQ97ByVcv86oAj9sOwMyTkMor8Bfx4IMm4YlWpj0TOhxYxpw7MCt
PUnwwsWhuFx5bWL2TU2xKdfl9g2nK2ZjlPCYAIRxjb4VBFjYT698jz2abA8coe4Yls1kQiVTaDke
5ferS3eMLvlom0uQiKAD1xLF9nXiPEwpvnr5kH2VefZr2PPf+rb2jRTx6GtxTRgz6HBJTQaiGSwG
RRgXDmCHNe5qkbn0yqUVHadnUEFevG7iVJ2jhWwIoy33dmf+fQCBxTIg0lemQ/BCatnX7GLSsQcB
QiuqDltj1D6Bhq/9X9jMUxZgtHJFB+Y0V/ZLof04bua0CSACQv1hdjTXpQTlH43JdxaPXryLK/rY
aTgcmDG6HHFGuGFCwxqz7ThxAnwxswN8PPWNPSuoLk6HLlyPMkXkql5psV9Fs7v/Jg+d5zmONBXc
Bu+6aut1k8wLooKYARmXui0VBCf7efWbxclVYq7gpR4o3iM5e5PG59KS88m1mnQH82acn3+IU2ap
B+5ooZmfKT/CzFkNH9ykWAuqyLJX8ObylwEMPeKQEjdbqB11dRtu8KJZ8IwEzNljDruA6buhjmQo
L2Z7NDa12K4nFjrknZDUVlFKvKbsAsjaMaDP6mMRYKyg5llwv8WwYWccz9e1hskwGSEqKRbGYiub
bsMQ9R5oVGUOTzOMN6xhyIshrALg4jNdf65q5+IucZd4sD4PcmyRfsviquyWjeRuHMFEarRL5THV
40NIcwlEjRa8y3aPQkBazkG2DkuNOwu0tuEFDw9rPCnRc6b7JP6+yOrNG3655VNOVZM0b3Qxc9EJ
r/h04WluT2QXjiz6Mo+ms4Sqy6OW1X1eNNG0fbjbNqBzVDt4apyQN8vasNVCFYs0gG38Fv+YMdh5
TGYj9FBX9lBZPrA6kYWEW71jzeYPaPVY/38to2fXDGcG9mwvVcZ56RN7PAhXkzEnsEa9HzY4SXog
d3YZWT3g/X8iihs2mQ4P+5WYgy48UebTJm90AKOuZsOEd8Kq5EwH6xXN9qJEi9H8KQpQ7ToayIUM
ULP/XcBUhfQByHN6KWlBhXSJ7aqXO8c3nAq0oVaeJmnv38h9jKr9CH5p0ZaE3I9zkh8Q6jzL0fmf
Vu6EBIye0z1WFTploctoDbBoOrZAoi1b3PHAnZ06rqw4Uh120CohSM3MNAD1ScLU/GfKZ1kZwnaP
ciZXzsATUJUxQ9weIMBbiopYryiZdFHViZP40bpgY4UEZ3kpD0B+PKm9EMlwjkRohHEJyHRm+VIB
iXcNhCxhJPpOpOMiY6FJ8HlJoWxQ4HxE6vr8ubBVTb4E4x9blfttJJFcAvWAP4Kt1UfJ3B9/4z3T
ub0dMhIGgOYOUnsshj41E5PEq723S6e1fq9NpKSPFHYallEsGXq3VuZAXZWy8CwiN1YUwlxjlmAZ
0HbSpDaVSPeDSwAGi+5TfnaQ0f8RfxBQGdOHmM6Q88MotGpLhATdO/+gLMzciNC43JbFGj0HOpqC
5QH+2zJyEzTDzB5G764U6QUBlYzQGi9oRldIt6bGpQtnDxOULdbOwlk6TzL5s8X+UM6aHEhHM7r3
2991PwLUscc7Z3bAW+GtNoWRVNhzsr4IATUpzRyEpCjQwgR24L0bIkUe2gsqpVq6O/HOru1+8S2N
rE05mtrfaRU9XPJ4jFS4yMFQkBJ+frNG/qtTTpcyUTPTZPcLFrABAzBPPww52FNiSWSql4E7aysi
fXDnvmhUh2JkkkH03PwmOjWuNKC36Kx6/SQgA3Qj8HLVzVBl05vmQ7MJq41CTbIOYH6GbtapwuQN
z8ApKQdZrRuckLqosvrHzxUroiCKGg60omHXMYkFfBCn9+rK8Ud1Mo28ds27WfxWkZSFjhVKuHh0
Xvvkysnuv3C2V5xGmkw7vyiTjQqs6KdUwBli0oPR2DriUzWHGctOlqElbLUnifI/vTlobobiki9/
Rz2KVSGcJKaxQTeox9RqiPj9zBNvdlaEQHyWGu6Ym6um1g5riwIPaKrLIyWgai3yrKJFbcvmEWlr
PRVcQNw3IB/2hmpPjD0XIxYL7unMSVcvUwhEGqsExkhMhryJJZDULdLasil5yCo0fg8PhaoF0e1p
hDos/g6OBlh8320qoTuN0zgTGeGb4rhKduo1STbEIQno6WdqTKPoH6ycQwGKnaEcfsMMFNIq/DGX
Kg2rEqAnyGxwuw2v+xQCgtlJCoeMa58yxj3mS249WaDWEvvQm3vI9R+qwINvNRJbjt03z06ljA/3
Rxab+rOw6ZRLrUwY4nNL/dSSlbteuJkuALyar7QbksJnRnn7xK2gM2AXtQpogRDxNotqSz64tTJf
7+OC1+eD9kxk3BgrF04aaFlAJsC7WYKXCDJdV7J09tejK1YVeViPDwBXosLpTTgsCPnakYarjtfj
C0n61uasgmfHEQlFvae9E7saAT84j2zp+/oC5lOcaguFVD7RMIBgCjI4gpMoGSgF6WM4MzsG22CL
t6h2Quopso+M+TVJwkxUw7axRifETcgS4bs3D5V0fJpR1I0EyZrEElaZYfOXRRC81r1nyGMqbBjY
iH/Fb7Ro8EV/GaQu0PUxD9O9RmutmgPp8YZT0GnOqpuMdD5FO1g5XayQRqogjSsOufKIIkl39cTR
ScWDqu2t3xcibGiRKGoY5dg+CQHipi6xcGkZt+gngEfb7j7T8dfthK5FnhgqFDqZ46VRebRCV9b2
/DJ588jAWkYucOU8HpOhFj4A7LSumRh6Xmp8AN6Y9kQGpnzOLHwt6YZunC7wryxaoyQLN6cClks6
DjorEcsU7tpInItF04nyIbj5EUwn2oA+Hm4s9YiX03obnJ0ImCRHqkk5V3Q3oKZKn6LhoFNEcABV
SZh4DsglhOxySBBBxa7sKIPcNBn/mphb6c7QcVsftaAYE0bwTbXhSy7UZmBpSwHmUoIB03pzfJhM
b4drcGuX0CfW/bU+YjW344JhSt0o+m/5z4IL5VYk/w8y2Sw79OMnNfq8bAsqr19geJ3FfITM3VqU
guqLfVxZYuDyC9jWD6EubCpjW3nu+1/s30WjzoljxJX/XKwnj+j6GFF9J4UMtVFCMhfVlfxFbZ0d
6052depYrWR+NgcTbD/fMEAd4PbyKxc47kBKc3MxiOfMh4h7+3FND86anLjN86gYpLQpuJ6nWevH
D3jNNqLNKxJL2g9/Tk5SHmPyFnn3/wbunCm9xbO5iJhN8iIFot5FR88MvK6wsbpKlO9KyZK1u/cm
3Fqh6x/JoHDhD5WhHmlbHJeH2NxUvbq6iDRkVIJ9VP8++NgDAot8hnEjNcosaTuotK534N0Afiue
LoPrXjPM6IHosXK6QoGzmgcL3v2qCo23zFm2y9BKy/x5vGfaRtJZvR+oGas2305Z6Kfd3/giC7/U
I9TK+AGM0Rm45klXLg0tH3T5TnbFgHLOIupfHlijSRGtzeGO66LeY8wQvGXPDEuURp+ASiGsSbI6
ENCBguUxRfwgdPJmrC8Svm1+7MQxgOo0fd0lnrxiZVYzz08Cc83nPrZxvgLFZJdswKWGhHbdb51s
lztDmwgK++1CRXvIYZE1hgCwXBvJwsHPfwvn5qMIU+t1yt86GdfrRI9vVrG9mJTo/1jQEa89dJgh
z3iQzecLri+Sf9HOcON3KvkgCk+2wNr9z7nR4eYPRhMAZug/xYSZPxJzNmSaaNDt2zSSwyaOXWHg
4z7Om401ksW4RwzKt1A9IWCHvjlLlRCK3gTuyZ2YxiGuU19D55eBqxHNUDFV10/uWBkDylsiaHGq
tmdxRDYnd8gA/oB2UwrtTb/B6Yef1BtUg775m113piZITaAAWvuJCUoSsiTlJWlNzf72AtgL5vU7
rQeue5rVta1ZBSCbg1PTl/7CYd20NC5/bgbYvE5IYI5T64TFWZpmgNm3lBIed0UzTqypTqHauAQN
U36RaAc9onj6WJXU+O0gOueVJdhUqsMRVTahtB/OC69qHtp8RAvCJQNPYI5CGu4GXxutyWIHYRll
vSdyJmXa6D9aheAmMMXhI3IoIw5aZe8yownfvTAIMAdA3fnDEwAX5L7mZYD0jQMcGya+JahTzozN
LDTz9LmG3QWPpoFaQwYX8hA1FgRJCIf531HfmuCsIMlog2tT9lbW5uVdvdXdkvpNIUD3iS25ofxp
oLe9zAu8N6CG/m8a+xHzP3zIy1b7+DKd/twGVeQWh0P6wFRcXWP4RrNgt9x2IQ0Gr0Nl8Ba5X5pk
3t7mJpqADvy74ErV7e6Qz6EvmJN00e8z3etpBYUms7Dtz9fW7nRbvPA11STPLc9/ItC/qN2cr1+E
Jk+UQiMblp/rFgSFHp5SIg4SghZc2GiOUr24oHLlY4rmf2Fnm36k841HaNKauQ1aikzXDiM0zRmt
lVqLknrRVQdodWE4rvKWch/+G0Wf/C7SMiTAhlAG6VH3wJJnekqNknq+hpeHjkbLieane/ZWBfZz
Zn5e8LdiYA5B7vfXAgHXMmvnsex8i6xicZXWeZOGmV8uVpS4/R7Ezj2PXC4dfqKoEGuXYjhTiJ1M
Z0MT64Mz5GA2OXA0cSuSDHmInCnDhOAwW8ZXh43ouuCyMAlDSlU3aBO48MdmvW3l4vno7CddHXMA
kDGZgSNlSom2S2gyj6nN8vANYiYxTjOp3T5EVNV3TNvLDTQa/lgnmMsqOdQgYF60+oZOBumHsD8m
6nm8COuhRIe4Qc9vXj1Ne5/Bkg43+EM6l2cESInnTvYbcAv4/eQH4zjiMu4n3BuH2i4RB6gGKZN+
6Yjmd7Nv8fTXBlzmzYP/4i+7Nh/lLI/ksPQKRUe6fpQl1e/dHS5OZTT7gm9flhdQ8wh6ttrGtpee
nkL+5duywpbqxeRppbmnC8fm6W8Rc2Dpj4nDvfQPnVOOvgGc9LrO3l145RAwSsE1hoJPZmZ4nK1/
lsDk9poTwcXA+2hXXw9BkZa1GVoNby61M1p5RhUArG6zYXED/ruAOxbASXwwjTCFWZzVy6HaCU7G
JIF22v2izWgMI2WnkJIhfcsEj3RA+3ZFEqedtaLQ7v2XF0heRwB5B+/djlg8PNwMR7Dy4UxRt5Ou
Vo5ICjNDTY9/x3SHOz6ZLOjVeR2tAtsH3ph39xhOcfFukkn6IAexYXIR4oW1SBp2WMRV+OdwQGC4
1cQYraR40I+iG/XSDYXwH5PjdBHm+nax/6xczmrVtS+Xga/B6UD7123wRO65pfkalN0JOUfYCm3B
GVE+q6Bv5CPdQLRHQjR6Ac7OaG+AeTU3pGoo6BxKfnRwnKFlnrx1u1P5mAX0gkYKultbwVSiksXz
VSE3tr6/Nu8ooSZBIPl882gyA3LHYni8gJzC1QIEWznDxR4qtoDMtmQByD3n25HFsDMRHEMbGM7m
auAEXCOSvLQjIYwj3FlglwfLuvZfJx5v9WmEgvtCZV/hMPwJYKSA+92CnA/i2V5IWMIA2j5GcRWn
/D1wLbE69IIbqUr72I3kod0xuflL7e73hCJIQaUyV8Jqm5Urxfp/tvsauNGTI4NqEh0HDWLEeI3a
9i+jud+nx0RRsHArVh0lFtY07pEGdBh9GY/IQ068olDVmv9SPqUjw6G2HMtDMU48s+4PU5/g75SJ
lnRjIrpxI9raKDWL+Ul98jWEsEtqp62/4LaBxerjB7vxPePK2xE4iSwqJ8CDkW8g9hDubnB/iN3a
pXcpTsQB06JdEba1ws1kdMgcple+k0R6lVEeu/840tukqPKOn/dm/G9Qa6Sgatl/DhmlC+Qtlc/i
ZsFG93J8QjrW08zIFupOkANa8BdGkHVg3jPqNoQxk8Rh1DeFFMdg1trY7q6FSxCNlq0YWcv/8Zmu
Qqb4lvF+up9L4QIjPSLseu3SKs0FJ5TmNWhMCf0ZcAqJeo++2nJ9DmpCrFfqoF+k3ANNUytcp/t7
WUnduxpgyZ66gl7NG7+35mexR2lu/NgQ9AztC94f2Ly0+oN2IiJvIJZRQ5QT2E2rSEZSZnESNzK5
czpYAikL1zzh3sL8nZb1rxe0UdodWkUK2NRObujRXT1A4NjEgT5Io8MFIRog9Gjk9hA+fT36EyxO
DithF88dCMHsyHmG+pdAQWuP7U1V5fX8pnnNXhG5BczDLMJ/Bz2264lknh5M5yHXtqx2Us4y0E3t
BufOwkGiLNSL/kNMAdqlefSs1waeg/hfFjqe+uEO1Uzm7xuwBdtVZirkODI4qwuWEbcOJGRiu0uV
3NT+J6gMLSCk7hdSL5KUNSE9VJmuzPN40zyfClkGQ9FTxo/BYe0OHN69vt/LJdFQh15nFX/ry1r5
gEkx4fCr9iLK/nAgz4Oo0U+VIND1MavCOdUIpaQnrXTS5EOODzkfvZeIXqUeek+D3ZOwvcmzpeY+
9dEzecbwq7pOpPsexkx3jLOosN0hnfyY/WYX/g+vLsew2PmZd+OipqvgI1mhb5l9/uIR2cKAYT2h
fEOijR7YIlAHEEiQ/Qh//2kc3dtewIGDLNDKxQQ+18mGClr1i4Dpd1a9l+zni0x42tEomlivunFJ
24YOkBWTief2tmJhTjxiZy5W54c9VIaY/HOwhdO0cIBYCbq66GlAHesPFXQzBf/NJbFqPu53RpZs
ppNF3qHfMCeP3+ZuW+qMRaDfb65nXpjKi047MIT01SgRAxMEi7V0raMcgBZ6i7Ztag2lnJp3lNAx
8T1SjhkaGxVp8geAXbwAWAqI+eH/lryqZKHRRCx6BY/ORYXP3k3HF1R0HmC3DYDSqIYFVjyql9+z
KvKwZvE/XWNAyhCahJmLHK6pgKiW4m6agbdtOKfqj9yBUJA6XiXrkyM7RgD/g8gIfaw8bPn/3Erz
XMNL9bqleDLasl2LsGpf3IGV0rYeK/uilbVW+V5udWhWHw/v2Cd95GlHI3t78gF2VRXeUy1CAt+J
G20qfW0vS5gtxm31utnsZsBEbpEqopm2mROZ7AU4Ritu7BaYaQv3dTha0swEe8nb/ADPjay+oKTC
Znhz61aX8ylzsEWeg8xucIctXP1tVM6Em3imFJSjTqk4gGY+fqab1XyI9HTkTK1lo0VO45qkKG7j
Qao4tA0LWHLOus4svN2EAUSK9zRglbOajlW8EjAEJbtOdvTid3/5S44kMAWDhPD7AQcezIgjP0wH
sRP+pywNKJ2J1hX3QJijW1sjNjwoELG5kAFhf3vvTgTYuIwhkE3aW7zCSOQNGgDjBjRPl/gp8oWi
KlRi9ohgikohp+M6tcWjEzkl3gKWzAkiVaga89pR+ahgKIj4adcX/IeiJsx+WIHjLeyRsaByeT1P
GcgYofoQfpTQhule8cPOs7YZ/LINszcqp67kO42Vb0Ayn9weDZpIAEbXwbaqD6xHCTZf1zeb+GRh
ufCyDvllF5wq0XS+TVxZwlrfymjFbVUVj7I/BaillS1lmc5CijHRaOJ9vcRU4jL5bmlIFECigqoh
Dla+y3BEYvUBBFudg97M8zjfcnHuJl6WZp/OrL860C1yKYs1+1eW1nMKtxtir0UC5VyuRYQnRmAY
F/YZug8hCa2rISw6sFtYOjAp1qbK7DR60zKlmYkqbKe3y5fdzj3D7KuO7kiXwvtKBoQlNxlDElmb
r36/CpZF+TX3t5IeUKSXgv1g0hKH9tMu4268Snj7D6tH70qvDHaVmOp0Ii0+XtvsZq61T+MRGs4b
CxgTFJEyyYXNOXyULNpnpoAQ4Tz26CDDJJtBnjLX8b5yCMB/JxANImlG6dOATqcfnUYcmAQn/IAu
6kpW/Zxb3ddXxc+rIGdMIbiltFGNvPmg/EgpKa9tObGJ/Bqy9yZvDetsm5FyJjMPycmQr2pVfxXP
G+OjvoyKP+kfqv/6NfPMHDERME9KB4zcABn9Dgc/tQwjlFNvwj+VBXtc+zFKrZekLcvRZHUd3c4B
GsMe6zPvG3r5lW/Bl384TK6gLeFUU28BEQh8oejkex71OmUwKZkWrxTKf16x00woJXABmvNX7pju
//z9tdVWgqoyd1zueB7GX5pSnlgoxQ83UPmUFOwF2kt9HpCzFDrlDA8vKfZV0xc5rhzym7i7U3Qa
45oreu8WFxHq3UpF/OIXfHqPD/NoQguq9OIp+AaflBe0Kb5sGWCI0iVch3f3Dzo5DFE/XAwKz77Y
Mikli2qMHF6W7RXRMHCnG7oJOim+8uKlSCWH55cw443Ep76oqkwds0QcOD67UR8GjF2TQMN+zAd4
C+I8cZglN9zWXp4zRrVPPpZzaNAA186POqQhpM4PsWkFvFC1Tj1YSW1JLPCU/VkvTqASJm9fGiQj
aARvMrPO1biBPQUN6f7/Bri/eeA8HNTi5EIPZL+RPaslT0cLes+2hOyjMkb5IHRNi24dtrxv1DdF
BZPVeQIJvKvLgvJTEvwrn2jo/zaJiIVVP0rt9VSdmjdN6CKKI+RPgW9ZGYRjpYJLozqqh7krymZ9
OCY4vBZ0g4u1QDXRNKJ4L4vPW73JMe5kOLEkF+S0Egqc/BT2sKWuMIGFGyvwZmMLR4BnglBP1dWG
U5Ekm361c9Uw3QYxdUCBWA1CnOzHvonrZNQOizeLFlNaF8pUvQTfeDmDet3dar7spTkKgoeY5dMp
krX0ASvqW7/EoODx5CIt1GpkCmqniy106akWlY6irP3mJZ2YKVfEUU77iSjvHFirJIMVvdngMAlL
MeMZNUV8FCwPrtVIhTQjfIjn9/lQU9+TSwsYnocOxyJqdFvPSSrlfImLSFm/Ha3YTjAjXCLWkaex
MAvAPB5BbZjiXQNIJUsS9xgxQ+mP2wQWF91QOoWEo9kdcH0avKzv2SUWpRAFO2aq6NybB+90m1bK
WUt97DaRqydO+NaMa4Zb6t3+N8wwjcQ+k/Bukjssx4DmuzxoaU+r855fUunRmaNCSCxKGyM0ccsP
7gREBqWkTJIJOEwJvJKog8+6m7b7Ko8/7CO3JZWMPUfL6L2ir71Oa/rleiK5dhGKaMaVSSeXIcTh
bBQaKj1z+/GvZphQzS91J5Jj9MtDBCzhq+Oa0tNfQDiZeSLsqsRb0zyui8BHmOwLZ7V0qrN7susm
6k5xDelLi1oWb3YrH12WbymXJhR3/1hyx0YjI7J7+k0lSszR3ywkS2/qNgpZonGRfQpjOks/rXCN
9DX8TI4M+/sCBIIFY8pI4e5ckuljwZg9L2uk3Iooyf4rtfEeorg3PanOSUqqfTwoV7VZgcFRgPfW
6sARA8cS+veOp4CUzCFady413QY36WA/NdM+X/qpNh8tscdUqVDQ04BaR6PSpep7UrXEuqb1+k/D
eCAU6VPj9isjyeyhp3Z1BqzCtdbVE3fqtDwT3No5GTDlFbytJkp5cAjjHpdZZhP16sf62D7971g3
Q/11PnvO/Qk1VcDuDzcKoqgT67T5pKJvkTHT8Qs9p3E8oL2IYeH1SFedvZWb0dG2sFT1T+HE/MH4
d+xvrWqKXe8f7T6byZaQ4vyNljTsV6jPNEaDe9I0p9vMnNeXlhv6utB4uHCwTGnHhpNSegHsSa6W
nQUS5cTXLmpekIADA5cXml/gkGr0Y9iXvglf7IwgLABYUP1+withXjTLmc3jItxN5ncH/4eWjUYg
N8Rftlt+OLZyDKccJJe3UQu5NVjE2pSX51WiL/wuJd/G3u3AZtLoY834LV6W5SZ3JW3KeTniL4SM
rOl/Qyg4TmlM4nv+CzFCBi1Zqm6XWDaRYlDy2Xc4irwdOMHuaKd6WPJnK67oK+T16h/CRJHel0Qy
tzp65x1YisBqz1Df4gkJJYOxtLAwcgH1khtHJZz1n3DNvwXvMbkgRfyyBw2+fcvN4yXk5ENfjcTu
qbiOKVPXbV0RJbCgfMjDyNifX6rKKx2DKgwwjvKqTYlT4U2aH44VKlHdWTHxM/sP7qE9I87pG8Ld
1DCfMnbGYAzwc3gPNvY/ky4oaMWIgU2EgiE8j+X/uVRfLYPLj7/HUSkcTCJSdVkf0qsdZP4s6N5f
uhV9Ml6buaxS4qyz92th7nLynZ4XjsXwbYNFUlSXf5yHiA9dw90ZsI2ee8Cw1dE/pLzPwVhUHjd4
5fNQ3i41NvgDM4mPW8H7yTEr8XgzcJ88jjAwb7it2XZGRIPkMdhDEM3BTw/yvcQPvICdrijH9ioS
KYaI8NzSJ/HWHxbiNlwSWYsq2lPIn96uD4LPUvu/vKecCPjgQPTcJT7rSO38G4IUZdZND3l+Hxqe
vlKV3dtO8OUeTn3eMPz/nvnwtlsapE9Ky7bvu89TD0WLxaDH8mIb2PK2qydeJFaLiKAEenpBr33M
i/QY0yGTFlXdKOoW4Ix4Tn59n+p8arr38jC8ANTuSRDhWxPso0JIhFmkOFPn4WCwFGoErEtKU4xY
1kB8zFFUfiSfeu5VXgPJ7Go1hHWppscNjoin47qIKtOQ8NMWe4vfM6wKV1K5+e34TuuEycufdJdC
nGNgT5c+UE4ZJIdSsP3iaxbtS97ULWb3RqHdZvXvtbwpyl6yqHjk+eOigD8SL2DnVvLpDdFiP9O4
sPdjqHzm+W4J3kRPh9ugfFrT7eD2qJvcVJcWPnP0dcLyinWVlYgY3VFZgddngsJkvWKoCMiIACme
oT20ibkMWh1n5Y/RULtZNqYkA26EX7LNyJKNHbntt/qlHVHHu5fnlwnr7w/mpVqVFKtnfWUD1AFj
B8q/FxRwhrpF1AvnYnqG8GNUFreFNXsx3AbAzKD5xRCnr8P+cWFI008HhHoReJPoIUQcAtlt16kg
6V8tTQj8ZrzrWja1kM9v60l32ZZGUciv2cVxu8FSGRXnoo88BlG0WmE87Ywl9KxhdXR7UaaA4c8n
uJlAHBFRID2AfT/GoAt+CCH0AgoJDO4FNQp6STq31yJial+KoPEXC6y0DR9WsvL60FW6Gsvm+mmZ
JPMELJDHh0UDGcvpGevZkkaysHBpOyaodQ9t8VcVQ5M6ahZCgmOi5GVJIDsqKcUFkqLAvG2bNZu4
ZRWy/sGeZBbcO9tZerSCl7f8ZWHFN4gZcXvgTRHZ6QzL8HdpNblr9O1xsx/5cVaDPe5Zj9s5OVAO
StpG0BboOLGgiEtJa3Ct+aVFXq2sa9O9ZrS0d2sfLs7+yH7OUFrmdiWpxwsDNph3YYwoUPxi6/YO
EjuqtRFPA7bnXyqcLw82AWn5eLorl9NcUk0KUgCbeEud9Q6BYb//LqU2OrTArhVfnY+x2iKi0ZGg
bJW2U3mmRLCgjxaisQ7RmW8JtzaCZ61vF/6YGaao6aY+NerLk4eH5vBq1Z5Jz2zCn5HpjV5bRfEp
sDIftd7hLVmwA868/wM1O5HwzzDIfeFakcP7yiPmpHb66v4as4X4Xjo89w2TH7ZkBsYgZgbUEl46
2jhYRmG/ZxeYdaZZx1AMlu5Lop/h2QECVLylVgLxuvUgeyeQnWTF5ZptjJ+7A7E+MZd708TmDj0K
gGNCJlVlifW4W9oQQB7oUxDExtleBktejY9qD/wuCaMGVDjtq3tbQfKV9cKWEmv54Q6bOBm5Kx8L
1Vr7seWynHnd0YrCRq+bpRJtjWxOZFMmrau+nw2nAI6LVJiz1hqJKxTqaAFcLEDTTlfGKAbl5waM
MqwmRIZuh83PW3UqyAusXIFpyZ+/k+g5Rasdyg8xeMGoGrvcvdKhwCuKMFqUWoL2QDDCsFAt6JUD
QPllSW4fmhnFAttEHj1PdY5XDN/KLaKfQfLc/MIhLFMzAFziXMdVdXhU7AIY+i/3Y8/1bxclRgX5
hz1S/RnOOEUR51i9assoT30Su8e7H+oVVV0dJ1P1BPnKlGLwMX1XtWq5JnPPkrYlwx/Wn59BNt5h
wj/4hDud0v5Q2y1N0mlHyM+wegswqE0d7RItk6RphaNr4LLkL7Wi4YMTedDyt0X9WNI9skSOOfjT
de2S+T5rq5K5onXsF7n2Ed4dXx7ovCuQPMuXbCDyOPISeJ8PARnurhaBMd6/f+CyEUsicEia4vGT
ktCfCp6Ll++mJ/8cJ2F+w/ew3xOE9zXsD3M7PQJmIs+Y6deEAh3gNAi+wADg91zBcXgjIuhx8N4u
3G+9SBWfFwST/cPRvCZzUAYTWwFmA9DDm73M88a6D1WIpSLAuiBNyhICy2iSSQ1vDlLAFa/Fu1T4
8JZBlrbpvVva418rHyGCOaEKGer03Sk8SOtzqJ/IIfnFwq6jeSqIgo/WTs71C1A7Y3zJlXC2ASzg
2YF6RPPC/omNiOuO7OhESA+Juy9ApmMYWB6WiXfVaPP5fFJGe7KdDp7N9ltBdxdjN3dZGIAjh207
TCwLQfVFL6Z3di/+Ve1z5KYmunuNow0wxnA+9OS9iQvcTyJQQOzPOLQrV36b0WPZqqV4/QKY8C1u
PmDxRhQGpZi52JHotpEslBIZjBGvsDCzPO/nNerYfU0lUIyeV/xstHaHAsxfIUsH0cKE3miaVaPl
RMbcdTea6hZAA3Mc7oGr9KwrqW+F1Yl7VdkEUbU3mmzCLG2xmCFFAEVxRzwo9lwbZbXKAmTOcYhS
6qGX2tlADYZJ0Hai2TFy/YJpuarKYCgYiqECDn1ktBG4wzFKK3V7ny63OceG3BiOMK8zTaJbD1uE
Mv5jHRCyvG6H5GwZfhXUIVbAKzz74yfi7wL+Csz1UwM+f3cI9VSQgcj29MouzNVspIIJCGh7xT4P
BqaJV0OqdiZ4eAlu/DcNLkorOAZ5EVE06+kk4dLxkrDZpsx37iu4VxVE8FI8oKfky8SXYwZlEI37
bXj6OVjlob13cwbQPH3e58PNaYnpdt1sEldNOz2CJr3ct4W+a54x8kMnccAjQUCifutzhhYHQipQ
kGWFG+r914jnh5o11XFnlXx6yLj8PXkbL1R23Tz9uZ7p0bVYuBgIzcXRsGLfYsvxuL3yIKBeeWlw
bKXYfnA2u5jifL7I3O3kuReOFqkOPi8DMTRIr5hzX5917fMo+lpDuTXLyH8OsY2Mv0tUTU8XvZDf
PHEgM5cR8yCtHXfsOqLkgwQGj3pWviOCYbza4dXHWAIXcrgO9IsOWLzlKGvKuGiKxP4s2t1MOhM6
bMPRcVNzCIDIF318zjqcyrHaSejJb6ZELsYMyDzYNcG4n42uf7xgHvkltr5ejj9y5Iqj3WFrINWV
5BJc1F+G/nj849iBBxFADcWRBcZZX3F2dbPTl7+/TGjXWDi/DbPxtUX0ZkGP926xoYgHz/ji1b1B
+IBQ1nw0b9epwiaIAqKXZsF9Ksfkcsbok+0gN9qrzbWrTv7XXVXrB1lnj4q0P3Kx7Qq42BaiJsKy
Z+59YINYeoIF0lC/jFrxxKWT0IAA3ckLnv5rBJ35MpvnIO33mLX18wU90XLjIB5I6rg3JCrk9VKg
//Ws1ZwyCGI8KBMYBCo05N1+cdnZiLRN1RYdWP73Ugx5lnQz4nLDwL3sqr5bJBtIXvKFLE+lf8bU
JWnMG653gOzePhqzw1tqyMFbTZpPJqytDeeFiiBWk3WZ/d/i3hl+oHxNByIPBst6TjaEz80mDrzP
Xij2ITpyyCn1NcPees5I1nBMzVJO8HGIFqCmMziNms6FuTPP6S6TLy1KiGq35gEE/aBF9Xq1MqC0
vY2iHYc3TAAZZbCFm3lczfflIr9Ted0l+Azlku4etfu4sSxBPSwqSiGH0fDijafeiyq9qjpOE+oK
ryQsezC7kcvGlciBqHBm7v4bsX/rShgZi/WLayl19MTPieRiyOB0h7Aiu6wMOi8/Zy8aO0pyL+8V
zeI5hVgAXo1BBzAy1PdlNtlWVUZRjK9bvbtVBz8gaQj/2VyTFH2sn9LUkRtC435jD0br3vrAoCRu
FicX3nbbDStQ6XBy1SrxsFERW1vUh/PZQQLQocN+kLz660I9QFoZD8XOFfew9vjTlZxSDgnLFDqv
SjV2fiyBSP6nWhkAYWTdwUv+rKDIsDbl2rd69VY0VqDozRH+rcaDxgga2D5trR+SkdVFRsQx5dAz
w3hqW9R4ueSYjk0mVAxxQTokI2gFB8AvSlc6PT/10RkpqS9CCj0t3+T7FcsUWq6idc/Goign7Hy1
B/iGG2nKMYU7c1UODhTO+jCmH/UX8K7d+Z2kqLZAsekoWUVsaw1NIGjOrX462G0L20y2oTL3DHgS
83cBXGBO86JHXTPPLuMyrbpNjwHMD9MHzjLBYE85ynVsNOhoqtJ5eZj/Xg2kfARhxhp4UMd0+Mrq
ob89Q6B8kiED8QkzNO5y/2Z4zaOKt2GVL1O1VrTeYd+LAmNpOBqn22Ns79VuMXyj97w2A7zqhTqZ
Yd7ro3vVhgRZ1O2Wgf06fM7XYu6wcF6RUrQ3a9hpZvVMPEixtDaPnh6byfi42NIUM4BUj009Ke/0
REP61wOvSm9yPOfYoKJFuHATN55WFwpi56mZyWwnIUURjYKo+1KPvehcD3DL4eVgr6yBnRlZuh/T
/OaRE/5J9I+S8MszsJSVUcFXycwjxucmdn3v17mZQ6Rj8XZZ7FJFw/f3hoUQt3qXSiygH7G//WO1
mnp9dWeBEZpysdk61+cDE9TvhJf8FB3ytw2+FD7ALO9+Oc7ekuVwH/LPuDQ707xG/wtcT9jBSZ1L
IQajz1Wnl68Nd6LCSCR6s/9CXOzU7yBP1iwaKjIqYkTWKFv2akwImBIl/DYee1ZHN5mwoRJ1tsPM
SCjOOQgd7P/huQxDHK+PLTmu085gACZnRhrwcII3afENTeS/kvIaB/tHy4sW5GdEbGM/vFBpMNF6
Peb7vLXpEJd9duHeWCKiIki9WUl4oVE+0xUsY0hGCinE+Whpm+ZwS9LA2Wic4YQTrTO39d09b6jg
JxdypPc6SIikNRi7VCQIudpfQE9WK6baosT7/OyS/CBIRtND/BwW3f+Kvp0FzyIS448h+u9TQ1wg
jiPS3d5r5jxtUZ2zoL8c258oLnl9Tw7vgpI4QVw5cXskZcnXfqU5/vFDcvrjtBXf+DCpT+AFPvDL
gb+wUwr2kV/bYeLxnRrRzC5RHToszZAkiSqww85YQgfi2RbZO5H/OnIRxz5irCmLnAN1EwOudGhl
kep7m3BgLz/f8QljH11Fb7mTRnFygn20eRkJIyH2DT6MClvftmVrlLincon8A4Qp63pI3nbNDhPr
2YGG8tlLEGjJ0ono8ebKosc4Ps0dvHj5IM0QVpjBAbi+JFgQZGqBATGUxtt4Lp4dNHrOpnVOccUU
t79IpglVXY2vQ9tZEXZ7cjZOwA/6YhkPGU5Pn/ZP52NP8jrhLLy6WkCmuMIqAfpMVETdjl33fvhG
rmretNxeCYzO6OJHmM4qNI91M1Fyjv0K2qXrF7jO33Mmltzy1fTDwEPs09yNen8ia4CcwZ38zj8I
OlbOf1NCJz3EMoS4IuFS0Zt5bV7a2UBlQkuh1HOWAmfxFU5uUHeg5646nr+almrtZK5aknbWhfzM
dOsIGafr4lwGGyB8a+tc0ovMpRqq9kB4CY3Hgo1WoCTjuyPthX55eE/xhvL79cZ1Uj8Zcmnu0V/X
wkDVxuV724uvodMjh9pLXH0MKAXqnp/zu+uiSWaXak2ZGstl5a4ffXxWH7hyRXS7qeTAasVoqeL2
2SAjkCFHSgvjoNE0LkhLOFTOdW3L2+mM2zQdzMa68YbpA/JgtQrlwwxXQCbwgVi0o/m4LY/YMQAI
TtHlS3/AKUNVlsFkqOAoRM5ek+cVlfrF9N1v5KDU1dGcR2U3Um8sDG+Pvn4rPWQy247UsCarsQRK
TXvon620335bccsjtS6z3ARJePcOBTUaKaMxyoZJji3epu38JbTx6r7LMCrOF+TJc8uqmIAAl4en
BO6EX4rqnL0lTKYe1CTykltbrJyLd7RBu92D47QxB9VNY1OM65lsLKUzs9I3Z/44dLKDukrYEQho
e5jQdE4po3MgRvcXgPiIcbXmvBPlj27rcCHCgVZ0F+LfgSdz1FNP+morFLGuR5r6hHevjeEdHZ6o
96anJVJ7gpnzI5upOF1HFSJHAhHwajw1l93QCfKSiZfaoZh1S8dS6rlrW8L16req7bEr4sPoagr4
vxMtZuvcpFDPynwFYSFUUcrxD9r+3XxCEIwxbs9Iqu2Y5lwUFSxrTPkv3tfmGfCZE7l4C2xmvLFl
rX0YXWVK+yeGqwtqD+ZM5pZEveQthdGtKUd31kWppjlgDodqwsgdLkXsuKWgTMq4Q0QN2+2gpTLV
Cdb9q1Vitrig2UhGEsnENormHQ9FZfv8iLPVyQflZQqCQNr9METrQsGSGbjcqpV3gyL0uBOyr6bT
N9cVxB5cieCkI4uQRjoxytjjnx1N5IvE17PIZ8dI6sKwAtiGwOMxYZkVMs1KqauJPKARZqRD44F+
X8wshborVRw+A55bXxn64mq6W1ah/SZhXs5x+3V+xUivum5d3GwjnddbxwzkWeLlWaRuPSbVy7iP
28IJYWud+QAYBGhNdyVfYvabfOiHrwDD2DxRbfTA2pU/KpLAaTKkiUO4Vvj3IzSWTZrGH+N6MGmO
+IoKt7oTHM9qWMT7y+XllA04tVtzJIGuHc4rJ0aLJjmt6l9qLpdsJ3FgWwo1aObF2rsov63BCTGO
LbMC4KMheqfr7sM2yElcPSj13n/Jb6ChtRNUnJbwAXD4nhNQGjOxx1foSBXa4ba3whY6L/z5D8E3
/UOGZX/jqYYpIKgI9/C/PNwqDKAAA5IUWgvwVnwlqyMDjNzVX+m9D2C1TvsmZkG433TBmzAgROmq
5aj8o4jmCRHnMj9bRFeJl2eo9V7THJurQCNHfQhP5qf1v/Eg8gZehLSCau+DCNw9ydR41b1UOj4c
gi8PoiRKDgH/ytHyQ2nQB1q+qL6K/EjrMzSbiBTobwTargg5PFMo/t49n9UdVUqyPyrUaKoarJTj
+Wpd6+RGeZhYnDN4V3Mou4xiKKZkMWyYfn5Xc1v7ljlDMt3+9IVdEfhmh16Anov6yKKofZFoIWmr
dgeIEOyHTYKS4V8Rh5hVM+9X0yrAvP/hoYOnXAySWcoB2ahGGsi16qYL6NnIBIA62Px1aruvlzNm
RVKMf2U01SfdX94lt8gTixtJJKXv2osypwGHGzMZUV9O6RYHG8bNppsQeHvJUfwLmeYQPt5oTIpF
KUlUFiawZppkagQF72sxGiKO9Hs3psASABSMkPSpi7Peadx4LmiCVtwuTSQ/mKychBnCLrz38bGo
URNCLpsyDe1wlo/gwGL/xWvSjl1mrdsJ5zmEmyhNX8PLaXcSjYI7olmVcUUgwTROvXEVNi4or1BT
tQFvEGZulZTA7YXnb11t2pT91xhZo+6+kLZFmWIfpF3q3V/81JmWObbY+69pksdqNkmqSoOatyQJ
1C0gIG3zg8+m4CerBqnXe4iWCrQBXYNHaBvGyZTJ1bZZCs36JekuO5k3GuXeTwqo2aTr1h02bMBJ
XVWeHVgpvi3xHFgSRg0rwdlTmywO6rJPE5uus+KKdzk3b/iuT8OKir6Ym9wjPZvbCMhIgXb2Gwgo
3TrB9ndnX1ZRzNpIV3vGlhCkzq8a0UXy7cvUhW7PhctGJWI5qwqKNgzWohkLZGHtpZLC0cSFhlEi
xe6BaU9NySaLMWpPtrhmawODyG9ZBe3qr3Q7MfqYT0kkBsZ2vBXkPz5N8htDhtB3D5CiX6sCIz4K
N89hoOH75Rub4Qi05rW9Ff8jCc35Psr+ytyRaVOS9+6wvSmE3hj42u3HSvsNgpRRA0Clb0QWs0/y
sXN1k66iSShZxUlDseGLDPliS4sDv27DQApeKejZxSpGp0jY1QHS1IswBjTf0H2DXQv2N9uDDZw9
UPub5Z9MULQqJ7ojY/fkoFqrGTnvpUvBfyG9w8MpPpqXw1Kwzy2QIZAzKJ0kjpWh0FPXUpi+Huci
D191rI58SjWRo5cB3RKMOGiTkaO5HYkd2m4SyS9+CPe/q/4fzeXvkdSzI90S+glgnOHQ86eC6aIq
zsN5R7h5EN2h5posyMKfXoPujqkvwO6yiUUFLaFhLIPbJZydEARXVRsVRjlf0zp13uOqzb+D3iCd
4AeRMAx2fOyW5SCJ+KKIsobx1lj+8RgBwgZPnq8h0ym2mK/fmIdA2rad4hWbK7dOdZCBzt8vMhXG
XOkjUtMCA36p/EFepz8ZJTQ4WpJip+s0NmDnsksJ5RqZk3yeHROWb7AKcl4YXPQBauODNHV/B41Z
lFUqyfOJjwY/v0F6MV8ZK5S2WiJ4KrdukeISUxPWsaoyQccY4qoxpcKcqbnk3vSjgddB4xTKB+2b
bBO4nPWRuZBf1kmnBHtKi6Pi2sD1wYwnX6UY6vCU+jrJye85XLAsEIG6cs+RUKgT/tNDFA4iHmbD
JJhqllALFxbVGA6hoZCasG+iaxhv7Dtl10BgJ28EMcqbt6bcPp1cdtl9xfx/0eysZrkvV2GXZq6y
fqy1QDbqM7j3/qarGRXB/BcnCI2dDoJXC77XuLuZBS1xJ2akwrdFN0OUwTlSvp6mw/J8hU2VlMW8
zWDtvGgA9uwFxZugoph2VGQF5bem52Gnw95t5hej3qi65Lco6LfegRqZKjiUYsxrbx5PNAMxEhlI
0+BLPPu/69jxu2DDyPk6yw93yZHAK34d0yOBIYKf10cZDnO77IrWY2G+ZkQZYGkrv/2pVijmMjAj
nF6fCK+la9IJyQSrrwEW/8KxMAdC0T2dy/JnDjq48OBJ1l99J7uBRMa0dL/33SytN+g36hq1w4qQ
qAZyUbiHv0AG8w9sPyaooq51fIuhRyQu8T3e5ZWhrfG3fubsSNanxx+etzxCSKOi8bdIm8W0Z510
6KSqy2otUFLsASTS7gd1125uhChR0j1sF026qr072jokB9hYbb49OcYoxASWiIIdSZcGWvOL99FV
nQVuLe06bb3hUG0WaA/CVhsLKfLWisCkKOPCCiJC5ii5m3iaxs9BsW5btYoDiW8B3VGRm/gMwUvL
t82PjTIuNdJE+1kqRb9KZ7Cw/MezbGOsATRY/Eeffo+GiobNBb+7gSIp9GS8Ri8GBSslR7GpRRkh
jKfQcGthC+xOZ+c9XwcqNK+N7Dg7hJqbA4SMoK6H6Fjq2IvNnCrpA8833TQrQu/MDPHQ+wEHuBFk
7WMEzQfwivtLPYY/zpTCr5/ICZ47u2Wu1N48eCM5ToUE+kTW2nWI9T/NADHY/jRp9Tcdb/iz5w8a
RNH6cyEd4D+DAD8sDaQf4vcaWY4rDYN+UpjTgEPoYpn/e3Laf7gDYWqd5NB/+yXaJLFaKij1mbN1
VWZwHLBCZ7fuj6xkpt2gY1bevbtX2tpgZ1cWRzXdXayA+/0bQ71uEaLXN7uHVaO4m/3OuBBW3eCA
bRLGx6ipp6vHYcynpkH11xgdTRAtpf8zfWPpr/jrSz80At8agE1KXxlTaL9kFE2NoHF+HFstp6pp
Y7u0g/c48PkcIQF3vqgUIZvBIXk5FLDxGxKcPTuVNHlqr7YmBncmeX5gnhU1dzmp13Q4tVrqt1/n
XQ24uQzk8TmPSZWQGRExmV1eMgdHfm5NOuFknEkDZAOjWrTkonWHBjkIleZn3yoGlEtowFqpwFoE
DvE0gen+vyRi63BBF8STAyjuXFDoLjSFAGTYoaCZYV1X1aOVBh5eYL5oXkAKjMsxfXsBnz/gUPdi
OQXjlC1mv3e6cLemj5o6KuD7ZOSs4gKtfug4Om9i3xZd38K740XkolVOcyH8whxr6KTKv5+mPYI3
fUme/nHPk2ft7pwhLb9Ko8XNRFLchf8OUHUXyvaJ6iy0IU7jahlnxVWRLcfDwZZodOQ7mdBay6DY
sDjd1d1fp2EABnPECWLtU5WtldhDj1d82j71l1P5RRX40HVAilRgkh5h6ZEs8z2Ykw8LR0K5p0R5
z5NcaJiwYOL31EceuRHfsH1H4dJcqWNBIe5vm6l1+pRTie2hPRCmSF3KmAbo55UeorehWl4Os49E
L3B/URFIHeeYNRk3QHD2fKVkF7BmJBvWPZ7zqQpsc/MKEF9I2Dy6bg8KEF1MLOwNBXmXfdgvq8kl
axhd98rYC/JEFFwp6e3c2kbnDkxj6W8J0DkTYhqB0lRDKVsKd1yt3wCI4nvmfgSktqlnUlOwpoPG
iefAsUXmW7jZzUGpTQPQ6V3uky+brAv+CQmfVGGzscTiZz9ZWmgYxePODDl3WrLP3Sg2gYMDLcqb
GsXPOCTnwemE6TLbLRxDeMJdZGYz9tta20L8b1js013nfP6quvhT918XP1liK8a9NjCeDoI5qSq/
f5IBfxg6wiH5XC+hiGtcKVnOZzr3IjcXFQxpXhAiJQ3AM02BzQnASFy5UVY8fhWFe8aPg0Y5EQX9
3pStZlLlTa6Rf/T9/EnWhTBHNpdEWM/wiJ2O2oeWs/IHDKYuANgrY/FWFQiE/PEbO/XaNny9cLPL
122hwbATiBenRXx72OPKhMnXgDlt80q03yVcxXq/VmfzohFj3lrG084ep1aDyr2/+rIh8rtxydS+
MVJjAdWBgSWeHSKlFGYnpwr4BROY0rcvmgek1fi3tkQ/ISFKTEkEVSiRmQ9BwyzfitJPoBvcQKoW
6v3VaxDJmInGYBLSIiU4EqufM+ScCc4zeSk/TfGXpKBAeVVVFQb7hQHW7Ojbc7Dh9+2sC0jfQ5qo
2E0sUROwHremhM8izOxPyzWSDu1HhVWf+Hg3n6or4UMRAlCwxU6r+T9eVJISiAQHBeMv5oldIsWr
aC6f8cjRWQiKMylHcCJOce+rRdycXnDD4u/PV9dsGXPbVQbc49u0XiAaj3EW1TWHuEITrgVvIVum
sA3jmcxGjzORj/uno2LBGC+9LpjOi+MMGbQGqgQPdxeyBA0jdTYCtd4Pc2ZNhCn4fuQ77Nvz79Te
6RHAyKyj0cdbRx2MxagkvLIkFu5o3tg5Wmv8j0HIS/6n1af6M7eVD7lG3HsZCe5BG1epMogQL+EU
qC0+82Cq7f+jwl98eA+j9XXV2DA69UkX+85aeqjAuXoM8duqkhMSw73uhCzPsaqqd3cIQXQUFPz+
J7JxW5YWlUrDrE7E13H1fDCkhsM1xEx1cKk9Jkj/xjshdiS65ULIKvJm0dEEjkLAjjadhRuDyuN1
hWy+JTESlMPdK1n314m83PoB65LH9iW9zpd/NEzJ1jhHFyy83Y2CpQQ/07iuqkjuR3u0wjfafXBX
HusU8kgoC9ZVRWVx65ahcdE5T/gEXn4KukrCej6mgZPNZeO+b6H8kl00/4O8be5SLLfUxiGnY+LX
zgPeoh46vGV/symYcmfasit6W6s5QpLTxHJPO3hOBhQ0LPrqtvyJWmH7+hCCGbti829F15if813x
RObItIKQ/0nxdRq5h+b3dvgBWXyOtFDrOVa3DMdi/5oWsheAxfxdRYF/k8kdtcFDghy2xS9KKm1J
4VSLJ9gtxdB3ePZXqoM2QGvld7MFkg6xyrpzeetUqQtjuSIdKd9EX3AcwqhP8gixgusoghHBF1bL
giyELEURD8O9xmUuELabGGsSc2xXHHRw9oPMaDeT/HvPOHTGKQ24aL4xUb9WH5qME+9vthwxQqxw
kE78vnZv0JB1xmMJB7qWXFcC9aL4OGhZC4WlJ57GQqdiSGW3MUz9nH0+M60fcX6yrWX5CLBF8dh4
gS71B+14LfInQDNZ+osM8OVx7ud/PRvX1+tJQCNjPhv08qM2fc48esc7eoVrpx9RVd8JhlbOqt5I
0Cdy1x1uWDYtJeARjPTVGj/FfV4q+Bnexka81hczr/t0VZBrO+FxpfuQW8ziCES1I9g3n+TMXhuN
8tJncE4Da+SFysxt3oSoRq1q2i7Gq/xFk4aF301Z2E1+wJ1xW3sbWmKHqvIJL5wdIWc1oqUMKZNH
LNj6NY2kgTwbt62zP6EJP08YAXLd9NqEJ6Wnl1YYGkOvTxOMspaQFzT2mwQlaJ02t+J1gKKM9H1M
8BrMXJDl+4FFT7BdkUwJKObFos8aKJkhC0p3gWZr+iUlhwH3jLTbHEdkko8SLbbXBnrzX2/mygwI
XwkWcWp1N0+J5+vc/ceL/9w3CHB9kyFKaYfebGV1fOwWm2jSVi0Euo7QrYZS3KHuzP/v+wYQ+kNO
4m/sS/jKUT2t20KCNI+8s5PqzEPZtSiq2QzBygPXnrAkBLYPgX8df9gv8acz6UGbU/WKcXX2x4NS
EaicNJ78Wfx6CuRBUzgdAxsnAPnHXrgJ2xTqqcMh7kTtHrt3N53E/kzdWNVkX68h/M97QGaB4RLG
Ql6t+SBKv5DV7XmarRP6iDlcJHCE4Veu+3oJzQINXuFwTaIso24GRg7VGkk5VjpNHlKQmlUzQPtn
UASPnf/k8cwgGWyGy44wvXjuzyY1Yvt7BQEe94jFIuCETrO9rn726iuc3xArjIj3lJ1kcVe4JkMe
n35fXM5H2DtV0S7v8HTU1DKOwXvS1/NPEl4yccx1Uu1Cc5quMZDrdhVweL0wjl+6me+vLG6tLzp+
7kRNsG8v2nML5Lh6iWW5CSjbY7ThnY6fLsZGOEIiA+oJR0lHCOHl6iGYJR0Y8e6IOZJksA3JAm0P
SuRibJVylKNFa/r261QeUlZMYti0cvtKzhxW1sCpXkCYV89hLpSZH1B6hBQnAhTlpjf0xTYCJ7E2
x8xAHhNZA6yV2qPDkOPgrCGR/QkShnXcBgfh7rNVS1yT00gKXT8pSB/LOt3eZJxQ/dCk6UrHjs3M
tCvF179emvLdl4PneKQ9HtwDJd7nHcU3dD/PhR55rt0+HV2FblqBVh+CIWO9B7qHgEUvm6OoqWL/
Sqq8cMufIrECeMI5EkkZclOv9SgB+QJ9pcBa6ZqjIAFABR8bejE9CoyMKS4nzGos7eMxvkgDGKAb
u26jf1RMT5XdFubrFm0aQADZjSIFohZ7oqRbPFD85rN6HIJhCEb0kr0wHULwkcmbQLFBa92yEtHX
oyAJUrkRovvR1vBeYhppTq9yRpwn/T6GDYG3X5XkWqMZxSVACfJhlu2VkeeQ/RLE5h0rwTwmCqO4
wiCgpm5sFogDF8QKx+gU7sNoDW8yBJUePV7flvK2viHqFyK/nbVYczRvw3POnbSz35+lfuQgz+5L
+0Y/McqcBaNqk3HFHL+kKIZ2Be24TSu/B40GaCBsMKIzRi0uc6pQdDf7H1XEIFAgI4Bl6wZYoU6V
HtclFa9gjrS+XLshgjaxnzCDFfjhVlOzHNxZY8gEenuyQ8PsqShIpS97R13fEIyWuF2iH0U/Re/f
TINUB/Q2XUnk0lmjsyu7uRmqIQ6IpCa3KDecyoNzm+tssFLRTv/9VQthEw8T6DMsuU8E4VskxEzQ
0HW8prXwyTUnQd4Up+0vn3ggzy1AhDlP79OWregv4F8ZJavqhOKy7t3uWzIgKSrw4wb3Z3r47a6s
oKXvcU/pjLycrvxoAA1iIroMlDlZ9q1z5Wvv3nb+XFGX53M+R+ZC2BKm8zOAqciTdo56A7U47uRX
D67D8fUhvqp6O6+x8g+ABl0DlZs6xpjSdaKxitYvcbTSBOPz9339Vuu5m37jZXv9KJcV8EBBWCZM
uLYEn4cMzNdyeU/fP8BnWbEggrBi1JXK4q7d4qEV0CwK4/fwLgMU8xNMMjzCbUpT5bhtWgejAbZo
OAhXQsVUCBf2JhpGKb8GqjGxGFYiHt5S0knA2rEgvEOPHJZADBGUSGhBgtmkfr6qWMaUSfj9ZaqP
PoPpbB8mT7Gx0+vcUIrdkMGo9CMJsIqwtan6VQtYJ/FajuvG9bqi1cGVL/i/S7MYcGNbxpNSjebw
xmL4JGFK3JvJnDuWS45Q4v4dcyfJcLZ5LYk1h/IFhtheiHy61wYyolDOQejv+gkx7/tOd1FhucVw
GfcnAhStVw5Vn3eW6tbYUS6vyfRGpSQSQ5sPqmdf7q1qdmTSLt6K00MpQSTyOPC7+BcBA5FWZ2/X
1pasQevaVNPhWmhBPz7kbv1uz9YTuceRQkdZPv0OIYib/TJhory/P11nleqUypjjv/6xcZ9ofr1s
WHlMHLoCHKKLvv9gpxTgbgI4IezZ4ffgIb8kcQPtM4KV6jRkHrCdh+WcZPbM/NDUb9cIonwkcRGi
e2FlLy7cOz7AdqOuDg62LLvmaUJIUPU894VCZfVXe7JUr4DEu5LGTRwxfL/zu5vfONJUgYYiydSe
FO1bKoaQ0xnmvjw/tE0/QlB1XgG4L+IjoepxI8R+ra+ubJZcyIhg/isRBdNlds9F7f7eNC7hQsXH
eYFyu24Q8HDaXkVOy4pdv8arqrC3xAtqRcBTl9IXTVHZkFIXC5BjeUHVIbHe/jlK+qMjfIorXEo3
cGUeKQfGQch0h05ECuR9y+iEgRK4c0ZPxe3910th0vNtus8/Dx9n9WbBHcfH2wh+2siC3FrmOi5l
y0ctDxa5ny9ELCbv9M8Codu6gpfE8iGsirtyNsQs5F7/GPFNgcquq3qKHjhE30AWssLuUz7osrRV
E5cA9lRgMo04Iv5MLrBTYjOca61QMbU4jtcMUpL/h3dzTHcg6amhrFNDp6tJLZM5hroJbR9bOJIl
7WmNMu92e8KKc8Xpw2oKcOwpypU29ySHA4IUzdZ2E+LF2YMc8LbEXF3LMD78c+/SaB8Hb8foHYhT
1B3kdpmoEbp/CzBHYE9QpAze1u15PIoK6niVSsv8O11P3Il6RPApsYr55eBQQ6YDlxf93Xt80R4P
0X6bJ8ShA/uCuR/j8yu/YDtMWrgLshZlN3TQrEZsBg73jjWIAkd1r/hr8W9Q4j/mjWFXvCf4jJaz
VEgPU4MFetST5WQejDMfWyWHNvCQjQlfUmlqiWgvowL+e/omBtMB91NX2rr62/jdV6p250aio1Eb
42Nx1awzAmAmha+zYSiriPLitB2ylApPjFEl9NHljuGaTHzlmM3OCP4k/WmuA6jLcmFzqXIg3Ew7
OSsMgdKlePRPO5wTpJQgAoFU1gZaUXCcDaN4umXI0l0uB7i1HFvTSGPZikhX92mpe99FHNrWKNWt
4ELo4BVPkRnJuJGg4KiQ1gJ3Zk5WIpyJfE3nlcypZV89VoWZU5wQ2+CG/pTL4RDzLzpJ0gE9IPMC
fBECZ6+47K2i7xRnlDsRwzNNq5eRv/kyCoZdUjnxESzB083wb2ByZEK14zuQFBi76PpUPJWm6mbd
jXJfyVqYV/2jhXuqMzQ3mUuE9q46a/737gYBzcmsxwlVv7Dn+d0UIci7V1VgzMIDUVNXj8Q6IxMh
UAKc/9/OF9Vo1WvJI2nK5P6AKHrhtAfvllABs88MntJjKfkyBy0SyMXl1uEazQ1UujAwK99Ebyd9
gwuYW12h4Q5hcvFPaxrAx9gcRWIveFYUem16ho1ZkQWxUCzUqiABc7N9YvGDWAgqhpUHjwbQMqJ8
NJUDnfZbHKF7vqz8xDfZnQBgk+yujvYbt4Y0J1LRr0TjSxb31IFXrb2jtgnknXhXpwj//7DvyYBv
RPOUsCDiuebaN2w+vDpn+kDMAbj0HM+CEzqYf9nc4H9P+CNnYveYu3PcnuupdPx+9NCMSSk7sDYF
T2tyraL9Dn3LLDKvX4uhwCzW0gesr8ooilHxNVf7rpvcQvoQf1mG8lqXUwL7Dxa+LdAnzfjOSlUu
ZH1B/kO4KowBqyJ1JRVVwTaZjLpTUlA3BILxVfKWruhZf6zS0/T3Mx+DxLk70oD+DPqtdqGXCOLJ
vko59BNIgjukUh6AJm4HkoIgM2dnFTiJatSyP5B+qfySCyZgOe6An8vF+YZlrf506+ZYG1XZV4Wb
biWsQXTMAOIo9Z4Im+MgCVAAI7FFfi9Q2Raet1Jn4EPrsrkYO03V2Wr+IGrdXlYfElCo3ibZTnDh
iqXOjMXAAbbBXYnKRUddoFh2xmWchv3xY2nd+hoYvoW7eozTKcOW/bTxYzkpG9PIAxPh+mj/pjLN
hkiaLOHsVaIVewVxzyJoEzQy7nEmRik3XAmugdKKFSEShd7i7yRbMO/oMxFv26H6FaXn5GlHOroB
T6tE5Twfw+namQj/1A1NHRPTtInzM6glfP5FvhdPWaLE59TsvYvokDGEqkqOKFR7VOBNO0v4IVzy
OOwHjBkzt3mgQtyTURoq7P3RTwYxxhu/9+UqF9JTWFQuTt9dmxJX76XJG3byO8dYB4ci5WTOb7UI
xuXRPELdYNeqgpTTMHhLZIgG17d8UUSFvYi0dV0lH1H4GCqm6z1VrSmWKdjuM4D2raNVLEZBGXFz
qLY2oywML3d2yDKBk0/QqxXlfBqQHMS/6TWzJ7KwONtW2mXGXMXicUi0hWODXAk7CEl8eW0WRaSU
qWICyoCKaXYi74RHRc/LUNj+14tMB4kqzWjdEsuIfor3gCrDqddAMTeVjloMvvNQF57MXl3MlWwD
M3h3ytSjLfm2Eai+OYsHumlYchXGZiBktcsWVkGs6RjPoFFLPSLjerwZMS57y1b7vtFdxhquagUR
4FxIwMFmUyJzuUfWlVMIpcqgk4HNUUhgHtY1NWP3gHc4YNRziHMnZuAt5Fpjcv4dpTjv7h79I5C+
sKRwrl8SpohT9sUfkFj+hs3UK3cmX3/TMWd3tNFO20icjqJK7UZz5GAdUteVhRCPdFuoSZeWvHOv
kLqrMNpovQVW2DXXOyjplgJq4Xm2Z5+Kjqs7x8z2fOKbxykH9E8bHQQUU+zsNMRUflweQizVNTn6
M/uUyiiSTWAzyDW1nj3joKmnyyOp35Ui+lDcSO4kYPGAibf6DFHhQBNGQEdru+ZAL4sohSW1b3Co
HKiuxH/QN6YVsGAFQHngtyub8gua9m4nZnrxJo5tEuE4gz1xKU+pCquRao4BjzBvt3mtYrHinQSn
V5BmWTCCWbHwEvZKrQm5YEUoMrtm/6yJ/8KbUWiSTLxBUvCRy+TWjCFZ3RulDL3ji4ULNd5bebXV
hZYq2skCmodcbsNpC2wp46fliMt5uXfNZl3x3GAjuVOAsaE0uUaPuB2i0obH1wGEoLEPXq13+M+b
fRxSF2Gy41U35lhln8QrPZh/LpFnzjHckL+i6VhFwCF5Ovk2wsYVKJqNullsXS0DrRR9fD5lLbHE
2dM81mLXbVbGHPX8rbbiDzDxDgcMNsJj+SdJLIzW+IzXpzN350iD2jkWnqHO7SGbFKl2LnHWgRA0
M6ZHlAR68/ppnm+vEKKFns9shKQBUuqCFcfLaibLouR9NgpbNcM6au8hu9qO6WK/OK7RTkgwAbfv
ak+ciUQKYDRL+UIMc0rJfWHMyYHMNOef2UsQgERBM8IzgHb7KOuYPMduCOdSrJgAICI+DJjETYkb
wEZj34TPVH1lqi2Pjip5GBt+1d/inXWvl0QS4JdD4zAq0OAIGIoWrtJeGyEyFv4BidJ1LIkMWV1M
GJjB99aoeIdF9oN27jwz48IlUFzEDadO4Om1sDBjD+R7//8m9xqbuEjIaxjbQoYQ/KhOjFDK7MI0
QQUzk7Sciu32yrK1sNHzq9cSMTnoJ4ypuLlJvd6Hz4EtnmnxPWN1XFEdLfmA+BVJW1IqYdK94fE6
YB+ZzWHqs9Iqttg/nkzDehoqOZIRfevbQnjGFp/AUXq7hS8NBcQ6zjgOT2QglRBATUoktGkSX/Ri
CXcQgZT5xgiYTtSqwhOer20cpJLaPEgsYLgJUclKb7om9NeMuNP9QUh5tkGeUXosHI3VlThNDOeV
9P71NlVjqK/D7nfk9sSn2V6AMiUMK5tS/STd/h5MiatPnpvjmVTntfCoOZiq0RuEGC/j8QkfXlya
XHgScmf0a2UkRHuMPntVFLXh5A8pHazKqLIJcFf2pGInHF/Kc2DABV4aAWJn/HPDIgw2LrRK0tJE
g+CM6nnag68TVSnyTJLfEQGiixW33TdOjeqprKOVImGzfTLrvGAT5dqhD0KCPQbUmytYHe50qev1
eYDAFsyKQdKiFi4A62/745tPvogvxvXSXuIo/z9U96hgihDMgzWbJus9MDXjH3fjofNZ9mWFZHcq
Y/EZvkQ1NG+jttGW3RndTZqUpm/p/Aru8jV8a6LiVmQLTbd66mjZRHRMmVe4cUZvaSBZL7GPlNNb
Mgdn+g4QXMTF/1d1kcJHglI60kIj+HM/qIWcrfEoQM6V6X8LxjPTT7NIxeQYbHHUhsuRvZhOSDHo
mvrNjaq+pdiQlIxJysA1UOjkrK74bfoAQvgrGwQhHhcmjgF+2cdqEUvRoL+wrL+buXKdR+e06v5A
Mj/IPtGjW7YpyDORrZnxkDA+3OiQl0UjbTSVNP3B0iNmGt9AziX+Ew+Zf1PvHbKv3KCHF6IpP8GY
CCzFxLw0nJWvEWa77N51WgWYV9w5OqtLfdUsmamxQUWAki8A6jvSTlR5kLM/gG2Dk8cPKGeLfIU1
rLZPRPeBM1po3rUF2K0P19dtYpKZSNcjjNmSQBYT61/eFp6tJw8XgdZw4DRF3bZZQlh2J/js7Mmh
xrrw6lo6ZCMT51xi4ZO36erN90FVx7y8AvunmGpLKSFHxtsDo1HFAi6kyC7iiJYRopawmqAsaUgi
d+tag5SwMFDSbVo33d3OMpPFOHkCfkwGd3MThP6OgLAdTTPfOdlzoKsvtskfoJ7Ief3px4fEp0NP
MrSrH+bekIjtJvPqs9JqkrcFmU/XcjXvzYmGcc7MiHGSpDSh5396t4iGs2w1+ccbZYbJdcdi0uPV
9tT2t0Jtx6AFWl5Xl9ad/BKsjAgdmM5s6lzoY7MTsGwSx/0sU6i8GH6GIn52rGNO9v9apH1eO+yC
WYqVlJIMl+AfewJQcEeljFEOw22MmySFBy38e6ws5dRHkacmc/XjZ+X3SGdnYWnUe17xzOjpd92e
wD8MziYTaLXZFklWbZetBmPB1TfFPDel2e96+b3ejvy/lbs5vXONdNtEVsuD2ogW9KKC6l5ShRCA
kGOO4akojkg7Gt4wQHTebGc8mkFeGkr8A7eVghPb27+GQTYk5ZU8/f1wg/O2aA1zd8MaC5kHAoTx
1m5e5hiASjsnjCw4JoY3KoMqMIUZA+GtyZ2T7lSBfQXSKsE4RHwwnEzNxDKiS79S+/WAOf/kIXFr
IQNy9635+WGUy1eDTZBUTpLJUVG58Bru3vvovQ/yQa0GPi5e1Lo8K1bAX2dMaOwkEkd2aNxvM7eF
bsXWUhRhKqrZeZ3JGpsBCAwjmok+kdeernwXaLWDk9BQaDBlJyxlAC45umjj9AFOQ2YV9zcsSpp3
1n4hBl8qI7uZDGfZYtjzbbC6nzsmBvd21JjxRXvr9FQd3iqIira9+sj8qEEwTsqsQkpnS03SP4DX
PT3zTyFtZzwKL0PicqY4COBTt+qa9RDUBCG1eIx++XmT70R7XqcwQ2wBmFnfjRxtcATXApWdhYbv
/2eE4SDr31ENb+U0TWfjN5imkWz9e9utiTIIJG6/+kb6dxK4fzvIZ1a4T4xdr1LLYKT6rFmiYc7K
2t8dKiuIKGdm42NPNKNwp+U2+x2pnOFY7rcrvQraOTXMIwSHP7XKzBPwwd/GPz4Ij4QETcYzijJ5
/Ah7zYGt348J9SDx9pL08PIdRz6950QYiL0LN1q1E0tJQg+KOFoUEsTODdX52+0nMTZxIm5yYn/P
VYsZP0JHY7PJ/kycNdoCeF3u5Hj0cAZluzxIank/js8xc4d+dGWS2UODU7aOgu6Hr6JBZ45dre3Z
6ne1t9+67J4fC6L8cRYvo2nz68uOw8PZCUEZWYK2V5uiejv5dlXU2PhiR+uMDaX6Igyds66VZH4s
2hyIWU3KrLH8L8fGvdAaX11yEnlipT6vTWy5GwxF4s7Id5iRho0ibiKuHHq0KudUeKiJaBbvmXbY
aUWqT7wInyjx3xlSVvBGh0Z+FK/nUhqxhLFjsoUdXTrJC+UoVynISw5qW+qQIRpqrrN6+mO3IzDz
KDaEzYHJ7stbFKjz/FR16pcTiUOgUtBw5P/tcHkqOYeDtvYZ/uMyGe6El8tgsU4qWq4AS88BR7v4
viC7O1kc4cbLot4Z8CpEM+l6AOs69ED9buDbuh8KoEEf7nnLJOO+M7bZbmjOePAVOyw2ZQRYsdgJ
GwetlI+S4BCyqDEJtX/rmFYRgelGTbx8d7Pi7rNN1vMPQaExnWhNNkqlbspHw63LmFTv1y8dxYKN
VHhrl7uhUJchcR9kj2R3dKtZH/GrAjOVepbfyqfgNRav2fZeBoz19WGYIFl3m5bqRLPUvj3bstLh
tShjIQfn4okox4yx1LEzcGGceOE4gCZhjY6MFNBY6SHBiEkJRgsP6a+CI8bJpeXwQCy4jhGLG4kp
4K9XzGS9nSOWrVCBtzY041UnJ4mY0ppQOlCJG19NsVN4ZtJBPBMBopJKTzs4I1a/U1BPmKmPGf5J
e2dwKFYu5n7pa3j2mZRn5x4WZULM4jPxy+L8e/qhU++LnzH2gFGKTbwwTaeipMQYTf9fRxPOsbnz
Tr+Wx3gAU2ngORHM0PjLNzS8/DuUjMZ9rSVnsAthXnKhP2dKw3cA34m9mhnR9L6clsfK/W7YPcU/
Be5CUfCx5FtZbPz63xxClM6tJ4wxka+68yd27wTvg4oPHACj13YBD9+J+Jj+8/RakYqA2uFjYIFE
8OB/2V5+Mvehbz56tlLj/gmsG4HXS+adQ4QbU9jwq2QyyjNW7UTUV2UdFE60P07yL/6yUgNERrvu
HLedg2z76hxt2VCXItodoMrCObHW+afg9WyBy4m5ZkY5jsX+w+P0A4sebEcGqTff5Di1zlnA5+Md
rb5YVj8O7k1V2pcOoHtzD+3NAo6ia+dn0qDBxzlSgYHYbOJFy0B3jBBZDc883XPVXmvpFvgcnGbb
x7ievMs9feSqCDEmv3hSRmLHh3klVN9p4O4tN3Q4qqkkSPD1HvLzWLVownrMnn06FqULgbcYof8/
PbZVC0NzWi2MS6NI41/fyEMehYfiaXIsJqaCLKWssRL9qCYX1ADxASAxmjkB4zl9KEnmamnNMLqB
4Hn9RAKBSF7ODHt0tD1PRLRxoylqbUM86dEv1aWrMlnIKkgYQONV6phtl80uVCwnCF+XtADF0/11
++eFIm9uCGHHE6A0Q8oeF0F85TSs7vXtfUnbrsAd4NbNX2QvgoMWBv9G1KhCSV4adGNa6GrmQ13d
Rc0ZUQaELdo7SWj3aOqElbTten5Ci93GCGZ1G3jnyCGfFZSk/WZP206WQk13l/NGRvuEeZBQ0nR3
KVIxL5B+XPhy1Ei/+mZHnmbyWQLlAiaI5dRG0UdRs3xcBuuqarxNHYyFvOigBG1nXBYvNLt091R4
4t6rUpGndnkTnkS8Dv8vB/gcfgj7WOzF+bwY/mgmymum68DUvhkXFLdtWAfQpB0n0itXDuD/wakD
a4OBcyyQBWCLR9ZiQE6T3aMOK7uZCEQzNQCRcksq1PeOYd1XhnRZksDOAwdd/12WuH8D73vHevIW
eY5WM7viR6HNzF+CHzgJY+VDXExUpx8Q1O3lyYl0KBNaqMM7P5YJBH52LaH3H6iMG8K1to4TeyPu
YgbIPzqDAz3DVdHH6/IMvd7DnUvBXiIcfQJfmpc7yCUPivEvIDiTeD0ZWk7iXwqi8gBOnhcLL3R8
OZ1opnq5SFQ61MceUrVwMDqJoqsDHvXoXz9yX0UgK61QvgSyjbc7qPeoXQHqCUNPrep/eHceVF4x
99Fwbx2rCJrTmFZItlcXnqnkNijVdTA7+ghFwTCLUz03rc1Q9HYhNbARQ6e1023zKX7X6O+drml+
uKCaQyo2ulcdEBiDS6rpCLydiB23P4MWrGI/za0qUHUOCF+ADOOlO9wCPzTfeb7wFOR5y4Ze+MH0
U4tS3aFp5ogGLTS2fEG343zXIRSsqaYnH+F14Re5j4JArSlHVeijJriPyYoEkDn/k+g0I2oBmixv
Ls6FibrtwtUrrk0cwQGcaTZ4AhopKOTPORjMD6O7fQ+gjP2U2WU+OkqtsBetmo/n89beKkcAZemN
eLsMBDNyTRsfSaVjKmCyLtA8XkfwkpNiiccOAuxTcXv9E1jtoZaGahDMALX0NK8gvb0CcJa3LnLB
3GXtbP8UOfJ086NuCP2wKVoTTFdpCd4IOcuLT3lWkalEZr5OJ9PTOMFBuCcXUmwEITlGHxfT7z/J
z03nRJiYPNhGmmPQ3ObrzKzhkYch07MpbVwsTauCRdZYh+hOG3C0UK3xBLpiYq44tV21ut/sHw8F
RvqyYFMUHTk5ylDXuHG7oayb/npDcbwGTymUuurhwwDBOU6nojdfsI9iewt/dst3E/3SToHYzHk7
iJmHZofgiD1C8bE6JAhFJwqa9dJgbQTBMbqygZo0YxAw1QdNmkUNjOXkdzF4jjoaRnwXZSmman3H
QOwO9pEddfvYVZCXRwwD6HHzkn4WO+IiZoqjC0NU6P2+wRuAPWOphnGAx6AwOuc85IVbiq76OqSP
Up7MdvSpcntnqSmR3PgSYRvOdfDfzYSNNUhqdTMCwtg7+hbC6NEt80IXyZUB1fXNIjp1m291yMEq
SO8xQoPg3FiTUkohl/a2p+91RI1sXkIo3hAUyW2zsNSArY4fEsyit1eQlzgGu+mPreOB5WxDkDek
FvRYu7uXVjNY1vWn8C5zyLR5C+bxyNBLNW3ADoXjPgO8Fb4JUKCLsO5tYB3T1a8rgXdTtf8WFvjR
Yor1Rybm/zx0J0Jce4FebCU2jI87Ztl0y30mFHtZkuoDm/HiTOLLXXWEXoRjheXweZuVLyMuSYH2
WxYkHXXhvpH6I2x8WuzlDW3rrtBEFwxqkj+OKizvitKwjp7t6mk3i+0Tmpjw/Wm5x7CVvz4WUPU/
IHwJzyk+D3B8C/Y5R7/JHXlGUEA4ikv8RoI/Bsu+/ab+Nic/dWRJ/LY95Uh88+GDKqZLuPmIdDNE
B+aFz+nAX+mVgIVAqPBoGrG/I2BoOqxD2bqSuXDlBnGx11ypUvUqMZaFIqokSXQWA/udhHdibK1j
m0IzS4I9Ou+xwYkTMjRVsGWRcLON22H/vgIs+TuIqVE1mljDbj5P4oBoXiBRb+H+AwlY9AKajWEr
y6ivxFLUdOySTxYPtIg/d0Szri753jSDZNCDJktUL/S/JGEtTeiWEQfP1k7F8vEj91sK2ZHQWOnc
pM0FrP7j9fpEiLsrSGkg+3yf+DKdM6w2mptwBi44O89PdWnQJ79e6bGq4Y1TFNxEIsIqNjCqsWhP
ZbWwRDZuLXa7b1Xt36ZlNCzYzn4pkQxTyPP3eLEa8FBtvsK9vgKgStwHEr15tRLzLMWWJuD+vbAA
+cbQByOcvtnmGFY21hgy3/s4caYhlNx2OH0GDb2RSdUoxQOQIadJjEywaMBemm3VrM4Ihpg5+YwJ
qtzG3Y8i5qvh/zTUloImWlDVyKsd6XJ/aKTw4aNdsHVtiJWz5L0s0kHOTfH+L2SU1vCeO+OFvzQS
hKBJOnFH/XP58QY5MEPpAr3t06hIz05sMLkDeacW7HOZj29q1eIri+HYc8pdpcJE15bp+iN+uWXT
uJg6o+Fddc7s6H9fNjD4fgtlhRTC+xHLFIxHat9+Y5QtQ37TMBqyyFt1GUK5t17kOvcBLxLWyhGE
0okQ/j/VrWgfz9xN0RdfbO4B58GKxJ0yqu2NLZTd1PNjuP+8YcVg7gKX+L7FAruBjmX4KfqGKdHk
lyobzDNRlQv3Wfvvp3gpiUUqAHvxR3yv1KHybJ6RGSR8cjJS17EuJO+pSq+jVCSfsRefoitWBB8v
ZkVBX8mE3vZTh/YI40e+/3WBERr4Fuf0meXdpmOyEfsmU8BVO69aOjhN7zkBp+FeTOxlhHebFlSF
MCLMnCPkRNI2PflklRrQM9BdgQXEnZQntSHf8/grv+X95UrceBq0r2Ig9IeH6SbgkUEG5MbX8ULl
lOeTKonWyFLNvtUSjZvXiZkkxw4Jxgpl9lbqdL0PpIgqR93wNXl5KozPHHf3AXEe4FWy7Gr/xewn
G16EWJ5MELQJlB03K+AwlRUxl5NUg+i0FGRAf3pagzVMtpuzV5HShIxutI9WiJjh8gd5oUSySw2Y
qpMwzpFRgfCWwdKj+Gx6NHFN0twE5Ea8uMTvYwxha6wq2Vp0JkpYCkc+Q+WyAs4vJBZiVc/ijXhE
khv777YV5knymFXHCXVUwVvJARQ4poQzuP/6Eb4gPtTkf3+dsaTQcEQ4jIoMCKindj985KDFv+6l
BaZv5NjG2AW7jAeC0NQnw8crgCTpas6fpFjFwPJYwVx1YfuQVhJHc1acDKBJ6La86fcuhC+w38Kq
juRe+trzPO9x4S8mEHrrqySOa6d5JEbn+01Rj8JLuJFiP19na0aFB7wfGLm4mvw22Coa3D7A57+E
6E3y+/yp1ZSe9ORpKo/B1PhH0BrWTppbU/Y6M3hJpMulHpCiRDMLCZxeiI3MzJVQAQr53n+NK/6U
Z+ROX2Z84D2gY6WfpeIjbsn4M+6UkEvRSuvB15MSYd+/KeAY4tP4qVFvtCgfyQWxG9HjcpNduWOd
WcoWori2ukiklyeU1L8MZzVq2icDBmnhpwpMRB0UFZz7I0wkW3hjm0yVEDCnaQDZ9XiBwIKWZCUK
LbAKOloD1LfvZDL0izK1jvSwHeWAg52zfAILqTBQTmZa71ETPRlUVBJv8Scx8dro2QHDyf8GvQzz
SXk2vTLWsCl4PTKnlqsWinvx8o9Tk4HX+PBu4ju23XElZavRLLDWfbdRCcUszvt3hjvSNdRva+u6
CbPV5NSfwE/gXM/IGYQmVncbeysdq+XYSSRSHiAD66v6dVLMzDOTyEgK2JutGajeu/0QSppFGH40
Pv1EpmC5yUUEjQXVbs9dZnd5pSB4yLzMUD7UNSIWYxS5ePwTR2M7t1cs5d8k3dJtM2MLlhWUC+lh
OBDLrxh3IT+9R70PIrCiTY6bgt+KtQOkv6WX7MbXArJiZ/QiYP1JBY1MbvqEGlSXvAy+BpEHNECm
D8GVq3l9JuMpp2XVmfJ9+zM/4pVPELmBC2hLhF+ehnPzbQ8BikjesyIH+7JZkW1czK0NtBYkvote
HkrZRyv53cTE+c00aYgFWR45IwDbuZTgXXR1k4dNRkYwjfCM2sv0NsvdHUyFMZMduC7HVqC4K0y3
+hAavn9BMzppkD1U9bQ26zUFWrZJter8M0GsbNo2KP92PPiB23e3NX+kUmjky67TeGH8je7LHxer
jujcyOp/lvz0LXwWoWrYrqiuNJJQBPEMJ0aQJi3agNEMftDsHX+X0FTYqP3SEYoUxfuJZfmXngbb
zF6PjwXzKnfOj3Q307lBpeVd9p6I9VsrbgqRX1PNVbKi2Cb7FGslXm+196t9fJunRi+eUiUq8AvF
dS7SvNfV9mBImIBSMhj5zatgKe4mHffV87jG7OdI7uz2TCvUIN0uYkCcfKURCg2otNkARQO9UxlI
FwHpLL5IxtIqpsL+g/eRDVSMuTxlzNhb0Sy9AaBsYnRMOtN/xhBRjlUlI+Qec6YtLVsiZi45vTHU
ViuCjfDRZEUjXzt5wJvn4L7oAJeScZ6nOi4eMm/ddQfhKgUUjbspMVlCoRalg1iP2MNgx1sGVO6R
PXUxeyC/jDcIw11qMeK72lxGPy8FOi1C7uNWQExkCOjf+2jDMi+o6mMVyCquqodVMj972oMuGDvw
HW1TVplMv0vHcTK4gArSIQvc/NpGaUFrkpoSUZHeLwueVfcaRJz3kCGk0Q5vTzyzKM2K78uLqQWM
HJH7kV3S2IJFdrB1q8QnaYgrl+cxmze6BLh6jJNJt+Y9zEqxsvQ3hR6GM6sM/T0KL6iE2qk9m8Ip
qbvehL2KlTu4C9D30zCseMoXZEBw2I6hTKqsQjef2LDDCaeqfAtVVdVyiJk9eu8VJJdOKSLQqFVY
fuhSa6B1Su+P2CbnhMsmqnkbxHT1QRt2HQK8oRHc5LgV9beJ8gzFQrTjw7xmKt7XPOV+ZlLn6gDj
EGcmn+sBVXmpaFZuEEYabikH0bMv5/ShOzF2mVoSBZ28Pid3aBYjce8QoDruNTYCVoWqubdJlTLV
rwb7L0F60UW9ui4Lm1hZjtZYK5KBA1mvAqrJ1R0otJQQrLtDyFaMjSZwy77iyUTBKY7WMucsPF6l
5GU14/mW6nOGGidUdNaYY9yTvrL5BTfIPPFIz/yqqAavhas3J+N9BDUFw9RnpVcljbXD6QrCraqD
98HD571hppgTFBrtP1rRyCG3vDd31zuZh74XeIek7KDwYlJzDb8dMBuywH/93s2/em4iHyBgQ0mF
SdCwG0TnFqYZNMde+M/+HYndPf+t9Nk9PRWxmG3hRoVhW9wMUsekYl+51s6VV2rM4t1unyWDIF6b
AAJqA8ENXLOX1B3P68FTteIjJwOBwEc2W96G+2kgG0kk5zXLii7jYKt6q0a5y0VU2DWZPJKl6FXJ
nmanBQSwqBh4+m221DrmG/V5Rsy0N+hImKA/49ng/oNnd5qQGHAWI6B+b+yS7ZTPICf2fVa505Gb
RsRWZbDhtZr9jKZjvuElKbLE8Qy6gSlEJ85XgVTdNdfEMHYrGKjMUQ/oz9wLOVcACLFA9cyi+4rN
sO5ak6V53nna5jYipAmGqvPSGBh3TUff+QiNgkTIDEcPty7iluIHiaO7As9BOMsckuIM2Bd0ALjL
ETJN6jT+EE2nUaaakjjbirxA3rFmZzfIsphAzhINmN59hDzRmS/tRP1nUr4EcDgNbV8Rb6DvE+SM
JgCKL04updCV3M/Ccg/oZnLvLYm//SDTOP6/gY7ze3/Knaf1MF7xZaPIT9aeYyLbSJMTJtZ23IGT
9ej177XVbCQ7DJXxaXZABXq4Uo+JlPPpWBHtSYE1zK/SBiMpb+szpBVfw4eWEIhfasP13ysW9JcN
DMlgFSKvpsVRLsac7W4VkJE4wsqW8o0c0lwrTpqx1RBwK4dt6KYh7krJ6wYQpnHRDlMduXHJdtBC
/20XtSHL2ULX2neBH77SqyIjAXdu0nxe1HTXcsZBnyl+a4+hcORR5AuTivcTE/bBtTvWFPanv0x0
zSRQrXd0hbPPM/FUu6yM2GhMtikSIh5qoUqKMsW/GmsbZ60CorvDUVciTqaM+uKiyX9Of5U9MbEX
OiK+OAk6tLvvyC4aNOI1JVj15N2p+TrtZSww3uDy33sBFdCXR5oRu9lYXXOmcm0wQ5icfxGmZqwx
JRjbnaSz7rG+SBlZuh0oj0ofbwk0C6xX+GizF34zfCdClwS4nvFJkR40oEVnJ90STGrshSmg3cU4
w0gkT3k5eR6CY6THj8DT6QUYmg2wz3jpdOhIfF7T0RDDls8uOKlccf607I2w1wd5Vv0GccoiuOQi
RZ07ZOlDLiAoftogBljPr6L30ZeOZCO0RgVgtCJIWVIfdltZR2+yYOTd+kyKCwQ8k/ZvTpdceDtV
IrCOhmjOEDfp+4a+C2H2benBK4Edo/4X85Te3UAir520GwfOHzjTd4uH4ReKwPjNmhvDH7dmwLr9
LRCtlLfmwkkrl1b93k7geno6Vw1Bx5MlbKsLA8clk6aU8qDTO4UWYRTfyJ0FaMXymIbMta4UNDM2
QYrC6bFbsRoy4CevpgptV78Zq5U7SXcxqtj+3L0HViSSffZb6MvnvZ2P9b8lzt6b6cS2MpdXIH4B
s9Nezp7cvD1ullKinY4LOHCVdsaEz4fzDWS4ONrz20K9qJZMDkS/4ji47rprus403JScjgtXFXyL
5efviIPcpQQdAy1kP/888zCkdWXtcIa6hMqbJFa/s94aRaGxE+wpQKHkEcrT/qt5nxAioER7ru1l
lhsJZdMSs9Y/SBbHzbTzcT0U32jEVLJC3C3tlFgQQb4E1qRAGDg2IrHxSxzqv9gHwSN/NfIqB9Uf
2DjuXoJ2vpZ2VE5XAdqo1twFGCtU0gHZKwzwSRWQjEIqQF4SAP+USmZmTbBlYCn4t4olBvl/ICtB
ht+Szk9AOVszGyx9oC60HeRTJ7SsJQKYTOdLVrNw8VWc0wviDSg0LCiHkx9v+lEhjGccoVAFOHe/
rWDN5o8FWFINLNEiN9VwDA+i2iJzssaruUci/UvGZX0CCpc1l/kU2elUSNkoS+9j54HFcCgV4SKQ
M9zjlHm3nH0eURkgeiKo2ZrwQ3RQbafuI08ofQZMOUA6fo1Xecfo7rO9QcB+qqvbAMPxhPuEXfwR
qryAd2P8RruPoJsiM8+91Sps8/tznqgYndb7A7J60EnxfGkKAC53nyvQDbD52Iu797kkcXZhjc9z
2YCXtFQJRc2MzOoSDw9RD/OQ8dtK/kQBgq5FHqdmvhHBBy4hKYj8InfhGcRg0BqsIhpkI+OSt1ij
ItfpKfTpMN8aSgkyxf3mRKfhLKd/1GcydK0xc0+OGJKUnGLytcGIhtwprUib9/JxQmLmwEQcxH3Q
L62eKBcEQACIbq3gNgBmIMurM2qDtnYfjwAVRLZAuatDk360DYtdcD80KDQEihuCqvIzOxU0B4JF
D6koFfJB4+OX3IMJ0PlLTxGw9ez+y6fMJTMb2Oquu/v274sAM0c1e3c3PvBZzI/c44okJdnAr6Xj
Us4jJ26qI5L4FLkMKebnau8K3vKpNZyqfWdShG/C415tywlgLgGAyIRWWpBoOV432WtxdH5/9Obr
8B4mXJ7igre7Bq3t/3Iej0CNgXRDS04uMViVujcjoqG5kR9Q+SNQAG3gnod7FtpLuejT9/VTAtAI
tMEPaLKpjDGUgXDKfRqc2BayQ/HZm1P0vNgSbQaqmtaBNWhnsYFJQHKLRQKpZ62A39IR/IeZzVj5
sEEP0FYstmRu2GrydhDLvd4HSeRwSejjl/DtSiHnO+HkRHhsJCKhj+DiX8As4ugl5RVEeP1iQxs3
Hd81GPvHz1Zoy9w5gqFLJiHKPP4B2sF4xEtlQfeyXlfCAwMhNbRzYYny4LFsYTFWj/xS3Xo/a5cV
cCaQ+uXAaJp62hI6rO7j+IuDXzm2ZK8onL0gIzFi24SYZ57YbynhFJKRVC+khXTNaJW1xNLD9eco
rjToPhsXXsbEyBMEX5VDGHz474n/qOBXueYfHrbuwRASkgpNdkFVOOaJqkIVL/zHip+KVKygwY8W
J8rUSZoPRZnWZBxddCAd+XJLkMGSGj0bhBUh+3XhRvpCP7aJNY/IDjdU4Q5vWu2y0WhGGF0QGP3m
LDJSAHoN7yWez9HwDGm9LroUqskOIwl71kKbf2WHkXTIeRLs3rkADRhKCIM2oiRL491WPqUlsCmA
XJZfAaPX09bDFese/zr84aPv+mC17MRfC5egE1OXQvkKAZGKAaxhpXkxQeKfAKQmindpA/2ocU3h
qlt8ricXAKVxwj6dGgC1BEMrswldazspLH2U6vSwCVwFRXqa0JfKFWX5B90yTUk7TVFxodzus2QZ
fewww2lj/yCIgzVUPdQ3Os3dbt8W5qc0t+djmtBBW/ZC5clNvXSjmUBhmiXBX5azx/y1Tden90r1
cUgrt6GKqoTmkYaMfli0FxHuw2PPSH9TdULeQXkjWtt/9h+UxFepilGeJStLoWHDr0k++xzbBJKL
ZwuGI2/w61jw3Taas/3Td4hDuWeLkeIO2irYYFKkKnW+ItYzdA1uxSVRIBgdb6XQG2qZuSOGYWYe
gWVuPCW0hdOP/5WaJzPieZeZe69tFmKPZUYA3OZa5KTHLPlifzlde2dCPfmli4vtwo8HVS1zKCx1
ZLFYTi4qypTEdzsSRgFaHvXMy2vpIOItirgkzL3RY6LOAxzUpaYZ7BGy/z13/XjB7utnswpm+R2F
lBTLdybgvPL0bZlcMdklRn+6VdBshH6GXu5fklO+2yEI37HIW8e/uveKJGSwU1Ly3lwMBPZmoQ8o
tpA0JpYgypnSNz4IJ/HVQhTkdLrWaFmDWI7AG/UeZEYLibwznv0t/yRyQZPGfoJEbCb1yjQOPHao
AoDrBM8ZShsFVY5RPlrmNrGrshvr70sehcmn8GGUmwAgZeZLYUO+4yIQOVrfhVAfzhkyn298DJjD
we3RiUllJsw9l0LyCQED8qgU1giEXiSQ0TFzLKH/BGEwqsd36RvWk4b+ggJZKDuRE/6YVifBlhSz
BXTSqKxVhp9XvL3UGNYNXjMfKumkBWGPr7FFpO9EzN0OliNAXMKMsnCqKou1b7p5xHaUHhOTiqaX
x0PHES92CEWRQxRiDUum4QtSdS7GsWnCo9UhKsezfuJ7YCdZTUelrIGaG8akBryj7h9N1MmkqEk5
TZmMLSYGi1m2WT8Q8Oo9lgq233xA1CZbTVv+UuFFQLGr0nAdardvXFcC+l/i/Wd7tIlyY+utoxl2
4CRSZeTrhNbNjjh5ygV4czi0/mt7o4epxF7LEiCzwLGgiRt1qbk6W6IXDpexXNgMt7XumNHa7g/z
Mvduf1Q43WwaNWqpxVxNbBtZjpoBgTPQXdcy0lqGpR1d6kZ99yzUOad3s3DDlFNfESM7MwLZGvpP
VOk37r1wsuxlfv5ChOMjtcw/T7R3OgYApqQzr1qiV9Es6z5lAo13YVh+edKsG1iWhm/cpi3mi5uz
WZluOQ/Nndun6f4uFqLTv3rkL9mC7z6YSRY4YNou76O7jvqf/Pw0gxmlIK29MQ9hG5adGvpyZTp0
g0bnbimUcIcEexZ4W83soby3CAxphpH/K5cAiaSo7kaVT+vTGLIPXWPGN9D++JPRwYBwNU6uA/4V
1rbfRS2W+Jnp5YVbeQThqyfj+jrnLnVCNnqHeB+WGWGTfjGNLkwIVBQwTc3hTCysK5e084DeiO0O
+/kDANqBuc/KYqf/yCDWi5Z5kB6Xvu7k8QHywMFSDx/R/GHK1knbRMpHD0HxIe/L5rly7aQ4PPne
ozC/YPPhYZWdRF38tOKHRGNXA6XKNGUIi/xo4mf9LY2pQFrR65xLzSge7olgh7YMeZI/YUji9IZc
ZSSGHPtk5jvf/4VndSSPxABm90swd3t5QDIiG5XXtBoIujVgqiwCRjJN/uzjsTMfh8WY0PGh6kNq
2rVk2F1ykeyZi4qqsNRJJ0maAf5S3ggDllEs7wSKbomT+Z+FFHtc/9OEFhlz+3+NmyhBcRWQxzu4
1CFHxLBsIP3oF3z1TwEfm4G0AfMFZNXBvsotX9urGsmvr7DSiaJUC/cPK4Ot7bUzFGAoeSiVhMxq
WPrxn5zdDHuyiLwyl36XKN8dkKQ6SEN4TH1aC9OSBhdXA5P/QKHNJczQg683ToZGvUI0O3EE+jOI
WHRU8eIIKfoZINBAEmzj31Q2cjmX9gSPJTSe1H0GdWAMOg33Bzr0Wn7UXBHzRqdwYmJx3edXd6Uo
kDGFKSnbEphC5TfWbNRFU6lnK2cCtJylqOBdA7eZJFvhOTQe8VjECagJRhX1GNqVe2JHDKBplrB1
W2Nkj+np2wAmnaSFK47vmFpDDJSzGyOKE/gbPp4827yzEdun+Gm66mwRuLu2lTgxBP7k6iVeyrnZ
kQ8YSRtBZiQHWoYo7fYdqliLojmWH9Im0W2OfAygxeBAh7LVcMYtx7PnafVGWSE3be6d2g2okrLW
B6pPkQ+8rHDW7MF62odFFEci+jIZP6U/mZ4ZV1uJLiI3ax8+wtwC/ykiCKOwGlZlFJBU4YDLrwpM
/g/ECGEaBBNY3nO8MUEs6mloG3ZUiqBMjPkJ2lgXGpMN7viT13ZMZGYDHBPNKOEyWiPbdnT7Ja40
jqglckdeIu5TvZkcI3d/IBiqOQn2JSXXsdIzw2rufxcLrQ6tfmEtmz+qPzcGAhKPOohBCWP9uh9M
I1aXz8SHZIAS79qgl38744wtCYpDeRIvLjWxYpKEzdhnATTxbnxTQwYucjUsNJcGlIOEpOJN3W+g
Pbd6/Q6do9RXvYWIVsG8NMnuj1gYsR1SCCV/YWghChqYj1Lf36iY25I+F2NEMgwvTECKpKYtivBa
ciH67efEPsVIgMwrCtCUKp13/67TUPedJZuPVNVRC+onaNiQSz3/viTdipRD4//9i8p4T4F/AbAg
y4QMrlCR6dv42X+VW0+gcN1RKKuQ0Yy0/bsBsu8vc12piyGtFZJGcl4sgOFM2WPHOQImkL7inqgQ
erVvtxrVKEhKjLEyANpgULYJFu8YBc9QqRn7KNr7JMf/yBxk2Cn76H2Xlf4SF3G/lkRxysnnmGqo
z6cgtZP+kQDOCCe6zLRcDaJdkVX402s6cwDTXAEcGXOTfXbUT1znxaIBrrel0n0as/0N5OkW2Fwk
P9wrM9J491hGA1iFitWYYsufSTKrSv0JKJbuayLbVyv/T6lNyTcZBrwMj3AjxJoVzrgQrSyXAOxw
U+RykvOD/ygwogYk7+l7DVm7vvPRQ6sKSTXoR1TR3y5aW30PVgJ4NgbCUb/OQjftnJv6DFaEkIDk
PqqOQ5dVHuX0cftJKgfuvcjUhIQfUcTqGAuJg8v5+A871k7vNGw4B/VPxxBRgF1N6Y21c0BSPg8i
ChYow7yn4Sh0g7QWZQ7+2vwrdRJ0b1ww1E56ZWiyz/BETSdtEOmev6n+DQyiXZau5KC8UxrjA9T5
Rny2m/K2cZxodR5oTf5HC4YkI6IIzDVyRqxH8CnNCT6v1Y1p3MRjdOuLWml6AsPkcKygTZcZWHOO
m6l8BBpClClF9YuINyujLmkQSVI3dBFJ2Cz8FMHQN2srDJju7UB4b50PVRKNozK9t/fASWS7qEx+
xYrh4oV8yHJObBJ4/fECBBVVIWnEiJW3dGzSQ36UH2nlf5AvcUcZVi9tKP1AhloWS88yBWx57o1t
o9l3wa/RtP9oaFh6/ZM248fOkPO8xiESs6VwnpTTfF9rOMDNvUPnSHrw7QlIdzUT99SVgIJ1HD5U
XnQ3Mhq/a91SM/H7ZJrhewU58ueB4z7VI2PW8cj+384oTY0rSdwgZStwIr5s2cNh4SYA9fnwNNBK
qns9ysWKXrAiDHR5RfgVOs+QfCOy+mPuOUXSCtd20Hyp/fpapP8afCl1bbjRA58jT1BVSVOGPK+6
cnrPQTEsfnQYPDPRfwx6tEWUJvVTbkwyMDIrnk5+ze7yGT65nCTDKUofkwRhExIxgS7rrn1/HxjJ
X6IMcq4N2kwz1eKH4eP3hXen83UusBBD/1AwFP9ef2guETpvszDlYv9/878TZUzeBuVRtgjGevit
U3ZIj0rZJ+KzXgsfnYlyiYaB++2xZld4LuTzAu0gulr2QYmtlb5pCrKzFa03EdmNrJAmfBNWDEua
F8us64HYNjJQGRN4/QbGpOi/TjIjT5J5/qWTe+8znZwDpr9Y1mbJm7J9zGUdtdj55QZcQj9syi0R
CADi8hfYEaveAqbzUXkG0njU6O/+PgYnFF7F/rnSR33QDYKLB19wKhwX4VNB6UtouA+qPlE7yOcd
KLv0+c7OGztWwJhSWj5cPg77kP2po8m5sQcfSP9QBKDfkNpSytZXyz2Fna+sDvIZdwBeT2oAfgX/
6WshXyWKpPgD7lZYFfuoOZV8MgCLpmxOyW1iOZPkoxYvdZUvsWirMB6ka9ZJEUsnUJpjroh/3qk8
GHGfd9bNn/9Fycecm95I89jTduLnHocGhG6ujyTYU5pXHd03uCGRcS1tP2A4wjDO9Tz7X2FfACD4
JbDuJRcXMA7M3sJbOHGgpKeOsqB90RUtz6k+fV9nlPM4PCNnVRdCywk3eR4jsA9zBZph8mfLGUMJ
5zkaw8ys6Q9cnP4s+zPLH9pHvcNaru3YfvYAB2WosxwTtvpFUk/wyP+Fh6JVfp/LK20CuwGNYrrS
lB5IGrklb47bCuFBmr0y5O7Gsv7XsPRk7eDZVPGD24s1JeZ1cJ/X0iLGfJDNyhyqjkH7Zueg4Y+B
G4c25LhhTLRsw++hHF8KGsA3IRu7UrMYTrw1Yx0cO4beDCsFWkcfmCWTop4OpwqJNAz3yMwYg1Zz
mqJjoC64m3vxKAYfKe/ednMQllPIHkY7SvIR29Hyhiy2hTcogCTzcdhMAmR2QKRDAXw5HiEzT3dl
Ju8w9HtOtyGaCi8HPSGy+rWBuRSOlq4+F2+E32kz2MdQJesCdyBx/kj1vZTf+VNrrZ6SGFkDLyZJ
rXl7Z24eNwLf4qYNv54rQkooisc3CG8gPiVzaPM1hifoeC+kujx5FfVLprq+k+O2ALG65/R3JSvG
ZWRPsvKGxhrn3f6Yz6y0gCGaJqbttbuI4HszdIKk0S2n0v6vqSFPOmKM5ywtpx/xYplW4QrbzfJC
0bYnNMu1+wnOtdQS9OnKz3RjHlR5yMBuswn8YL8KtMSoKm3WRpE6kRJFDV0J+Lf6CHkGQHp4ppM8
P3r33/7g5paSlK9eC5OQYhBW/e13J0Mrv2Jbq+az7HJ/qoeXjIgeUdkLiOCX1IJmT6z0OQFPN64w
FNbima6Icoy5WXQzzo9tZ5uhE19kCVe1OULHkSycu5HutAv0L3JhalN3HxmdmiDe673Axfy6k46Q
aReH9/q1QYXIJ4jw2lQy7lWC+V2LSggQm8nJ1GIMKGCnBqESm7f6/pLKZtnnBDb8VUM37kt1uGkt
f4bLKWD2CEJ7cL9cZj9Y86PYV8HYJUGl0WwRpp7tKuhgjwBk1XisrWlLo4toVr5Y7hTNO1Xu9vcM
nSGNQ35ZJNCjSfP39BwV8jWNIeAhmc+yDPDxjfwS0yEO1qGEkpDbOKsrfe7UguxND7rm4Ot7aDOK
tLaoIq9QBXIcrX9XXP1t6VcWxikiWZgh2ToPr0nrRPmRuRflgtihYkzgZX/YWEtM+xkzVKMy1CUy
mUIVD0FECSmq3tDkRqJIvUmTVmhZwmTuDzF56D4wL40M3ciJad5K1oqc6gWcXWmHBhUfBkPfCtIy
uhFI2f5hOa0Rp3ViK7P9rZWXUebGZg+5R6dqBVDW5hhCENLecYENnllDO96IyboD/mGPAxcBdrX2
B8rhWyspGswsFINfgNRfzblKEP0Com/fQOp2EBefz+EKd9F/F51wJ6x4Buk0AhqAIU5/yDOII6QA
9iqL8GnUvGTmJtw0Up+Yzu+sgu4eEcnX7nIVhIIxhH2KK4U7luNTKCYw+a3CC7tp+4YUox3jzEdU
jEAi4P6qpXhr5iTwqIyizkvX+hNDYt2ddcjpiFMZ8S4Uqd3idbUevFw9p3GNmdIGL0k2+WywZuU8
xYyhu2rHwfndRia00GdzKTffSGP7rmI1ad5oG8TRVH8PyyEG1U1HzD9E6O5N0xlNI6J+xVamd/J0
aM2m4DMszzoQQbx+a75VH8KNe7v7zGAt6kqATb+D+45CDsiOYsP5gpB+ja5b2soSq6Wpedih/lBA
w4VoxhHcIuXW65aegEspFhyJC54N1cQW2i4D2eWXHHD/rkyZHBSlZF3Btdzife5i2zEGRa7JaTCQ
kq1+qP+d34tBI8jiQiNqsH8nSuVGNue6Nhm/3pEzk26CsuKzKF/2S29iVCN/nA1EX0Q3AeyL6qkt
DY8wofVWnQdVKMuEsar4vCokm1XI9+3dlQkMdG8hNRT83yKVYrmA1rSxscWUr6+CZz7y0DVf+1Wh
yjZ5SVyHd/NQ3MvsZD1duDpa61MgpaX67pCzNY1B/0x3WRSTtESk9GsWw4/jmpf5TptSZAAQCqqi
2HAu5l3+XD6lhw3eXKpAE9WVcnbre7jiiWDDHo3gkNiJo801njYUtFM+B6VPRaHUZkrDF1PHwfJ+
jGdJsxBpJmiu9AUh/PFS+eqa4l/RXk+SXmqZP453tMCllANuC3lQHC4rTR0tvJlmIVw3vNU2iEI3
FfvrtARA/3YeNzuCgwLIUrkD6rPsPCTUDY79ZChDmyaR/y388pSPfAwPdJQgNwJUcEX+u3H6vu5g
gRgI/8yoteqPaAKwOgVzcAegAf+mhj5HN1BVI+qyJYDfc1QWxxa1u4X6uNFvi02n1MI+r5DCKi+D
qa+7eYNTfcyd08uv7wxuU+fBk0ipVlIN4QCI+rqPv6uBzIPj3k3KCWqwyxnDz2GmVzQ/eKwdVWD/
fhUxc3oztVh4vJVPuJsonzYQI2MxaMdSCm0yQFExrqT8moHJDRUK+IjmOGsDi4YAlWbj2myUfcBw
/spqcV2Ypw1X5ImwRX5GYgIj+3DnjaxwxQ+L9F/6yCbFO1Fq+oDqT9+SXKss822IO3OvcC2HTc5m
+8OHCbfRX1y2VT1qiL6g0hiDfb0iKVNe6OhL0PoObuOiX4nSc+6vBkYfIFS+7m7Y6ZY3l01rWEdF
4NWuacdxwNlCwmcj/N9njPf/5WubrHLBVh1+V3k1mi7205stWLONxY2lPYdZewMtDib7K4zTS03L
HtZQVXCFosKbvRd+yALYc+nTFvcd8ZGfnbj+/+oNdypKUacC+qWoiPFV3IF3PPW6E4/z/gnR/omf
kfW0Mr/hJV1G0kuu4SZMIeEpma4rWfRGCwz44XO2oA6oVMa09f5E6qQxTmLKnlf0DzLB2xXmbGml
HkjA4tE2JuMTlIbUHvNdWnWINO+5XlbQsY2okMoX1LJgpGdMNlzcdI7wYu0KZLDB8ToSmool9Bj3
KWPW7r2bUe190A4qz8N/PtmVtxdetovjTrmATVYjComSFyI1JJm81FHAqN0IMWCRn5pTJLIOIEN2
16cAAmm2WH4gC4N5g9XR7MqyVTV5Io2rxVg13rD/BLACjQuYHlfnv9FyDHs9pcLABcq+XDED69eB
xvjFdgGi0VYfOcbbYCkPBgWpTCehrhYf37eS48Bu6VXRAqdepq3YXMrImxWBqKW4tL35uafYiVrd
KwS9UuE4udG6RWc22lczNScuam/pLbkB5hKzGENE2MtUSV4mCoZLaYOB6sd3ZyN03C+JCegSJWu5
sR3fEhqF2e0jsvNQIqlfdQvRXmIj1YOsIMdBse8w2ZIWVB9ShKRsQd1NGY0rMwNGYPNBKILo2aKL
XOT7AHc/5g9XOfayBE76w+Ssx2Yj6sebqjEJ3QRKuMZ0uDe2B3NyIFLBqINIPVkotI6Ka+3Pe6u3
vIUtj2n6nCiK0JKZIcwO38y1Omk6Fxu3xADc2Js7ebVm6QmbIW21rhQXERl6pIYGvurf88O5vKgS
ghLgIfAXYCq6zr3B/v7iuXZtNxTqw/sSP+X2406HAmFUJa1QuGQbruOLfyFjipThmfDMYI2ADyja
cqIO7qy17IcS15kpMAXUp/MJR+veOhnchYA9liTOJ8iuO2gPiMRZyoE5yfxerebE7KHXdHRXvmYR
kmhLfQEBRLqyp58jy0wyffYKDiDEZIrW1qDPyHyQJvLNdWqct5bCIugN7AAIAqp2bkmRaQ2lyKAN
7qcBF6prdDn8Oq/I1qnDTxU5EprE4UhIGeF+OGfRWj6hDghzPwRyFUErbLQfiUA/NEM3jX1D0/m/
FuickLv4VWXBLTi9D4gWWxQR2eNrp87Hgp98Y2eEJYh6RNTmzWJqjQMw9qTfVGHw6xqE6T/WQ3nx
C/l4cKrVKr6yGYqMwOXG1JFhglZA5GEC3RGaOG1dYgUkWA1dhWpJiXlXa8vU7oZJTOKR5EroEPXJ
RTF9RPKiZ8pEJpqIvLok8IT9xxcZd0HitnAgHkmnU7E5AHZ5BKRMVm9AYBYOLE2B/1s6KN0itR/e
HZEWh2OupWg4bJH+44ZbF3K4EgJHJnotGUVrhkXHNaG7NvCeT9GXKUEFRJuGyDXSyS9bFOFns/4m
rkOQ9mycc0SlF3HUOi2oq6E7ri1zV55FFVRs6a/eQVS0taaVDLHcgF5+CtjlV5LtAotxyUWrI8im
CscRwbLSpGeiQDcYIpnfmIp2MMFzE2fSAkS4q3DB/4WA9yx5zY2DvajKiKnxdMZmXiXshz6KCJqq
E1FCtYNuR19QYfTGlknQj7ANCOs87MxM4Nvca5+dYHgb943dJGDOpEP32JsMp9rp4Q0lVnytjOfM
fmqVRTWX74pJvVD0+DDBjck5odVcX+wyiAyu/WZFAwhMkCIu4Fav/mv+dMsKTlZx1Te2KJr04zDi
9MX5fbwgo0myllpBRUjGc/+BZCld2GH1B1hVgoJvopvViSxr3dIUa997zvTXizEFgjyMMLYsNoMB
jlCru79UIx1xAnMpVPcDaY/KZwPxjcAaLavf2rurk+92mzH/wY/4zlEYVESx4aSif6utnCIgN0Sy
mOKVxcTxzwcDgfvruV2wkc9HtplqxEmy4QYyA1uuuJfX6mqYMjWByLVDzjC78r+56a9UO53DHujJ
v79gT9qkC2Y0loNqgcyJeZOJD4JQeuK0YOP1ngd6yjByf2yOaQpZmQ2ymMEMP6hh5FPH36DmXaM+
tU6+WweC+8C3tEME9fCYBpp3UsT39o7CkX9npxpozWGamJ1QhWcsYocH0/Cp46YsnUZpepUPolbG
rrE32DHFrcmxxEf/3REllPyB7wqbtWagugtmdY8lW5NeUaZKZURZEF4vjzUFoSyeWHtB2sADqpJX
q8Q5DiyPYl/qatJTKikb/a+x1+M/7q68c1NH3zpZ/MDyYCYkp51P1QDfLCeFsDyUzNyOk5iC+2ay
Jb0wF92NF2HCAcdwXNaSftIaBJJjJsf6scUJv3xTgZ/a99TEk5RvwLd5e1y+bwbpvX1g10qv7SLB
wU6Nb7DQROfqz8KbjB2rBCi1OT2A8oQ/rhqv6Z2ume5NnDvlHpJ2mnAka77XRxFlS8YFJgXpeHKO
o/188pRZ4/6UhhSs2LYoIxDY2HI5148rAaM44zAKeWd54PGGV4hER4rp6tZ7F2s1JrmHQoVQFWQw
/TOtm55cUrxv+L4sWEZmjn4T7y1X3ast0TLjDgpM1sHG2DVObRFwzzHY3K1Oh/zJGLkOhsIn3OQC
CCjKEeKsvCsn56PLcskXEIlzNHNVGz4h1nSpRDYSZhukWrAttYEznBvF3UZ4XDKxvbnDOm1RRz15
R5ZSo+iLDtRz46sdkksSbC3psgTrkdStroFPAmb9yqBWaEBidqFM1lJRF8MNU/Q1Evh5GFrTW6bm
QiwS9iwK7w2BSuNWUNM2iFYZwZ/MVcej1t05sCKqBIPoGvqP3tXlSR2HQOFneqdodo8BcgR/7YnZ
bw1WCcMRSEwhRJCuuFpyrqODV7PpbwPQ+uUPOLdn7/LA8FzbDGLSIpf9wQ9vuBhUOH7gnBsfB9hw
IjaHpA3ocjsUIFKQkj8HsOA7uU+/TJs7HX0PXqwCvW/PMTuxlnLz0or1MlpYW2RfD6fznPLaWeLu
fBbTxrqIv73EN993y+n2yBKLZ2K09v/uGfcZTORtlwBiX6Ehcspdj3RmKCCY1riUubBISTpPd1oU
tCnceFmWTdleQDR5tYlfELMSglEZ/JVQGiO1QJ2EQyw+yD/c+TiRiyGI55PO9rVq/QMX5Aj1Mjco
WpvLp5uMrHRdzoD7w9lPU4JseMBuUXENaEKlQs5xkN2UTPu0RwK+/kg/UG6enEyrmLjGiJvEzUYm
XoUemfkh12J3IXxE4prhdo23ySfkUas8NPw8CMIb+IKtHmfov3eV/uzMMzHEmXTCE3tm3IXRxhqs
KhhN9vcKuUxzfvebZVwjdueZFFXIZy9skToiCvpR7NYyUa7uzYmCkCoySGvIlvy/Mq1B8eO3coCc
bNuy/g/tSzQAdzdXo2XTppFH20mU2lpmZwkidoDTazio5cm/YYS7XL6/tEOdOo81iXEzsv0FnJFO
MoJoOa+eVsI5zbTNKq4RDZiCw0fjbJBqry1Q6P22YG/2WIRa7ZGfLiV2Rxrme06H63kZo4IPrr5e
D8fnaOYT9i0l2Og6jGaDmMaWxeJbWM1xyQgzl82fCYR/3a92uAc6fsETZUbIkcZrXYbPMM6rupTw
PkMc4LiG4UPcARN5sOOLN3Ul5JWyOcn0qN58uuXAGgRQGxZPDWqkej59O32i5+Df8BY7u03v5ud/
roIfFWwNVNjA3fFNZioD4RrXY6H/VCm9wsXevtqGM36zPAd/trow42pQv6AsJDna57Y/T4pJhc/i
DYbf8CQB8zjiGW9uZRGQzu1OI0JuFEU7tvcqFKjK7F67ZCzG2owkykrWoIBMxvQizw7HIxzLVLUo
BQiVRKZ9xT0V2wYg5TZ4RJrtFBJc9HJDSiUYmTh6MLFbQmP5HPEvAoHIJOfvVMUY+SNnQKCiPTXd
Wb4B7ADqng/Zz3nY8BwCg9I6AntBIAY1tN+f2HpIzY4UISn3iwrUXJilKUoKIJH3nkSHHcMuLTOf
krKx8Pvn1d0+joeaLkW/Qg5j9Z98dth94HDu2ee+T5h+zLn8yXw4T0JnDy5TmBlJ9bvR3LQuT8oj
u+9OCVOhczWMjJMCxj9QSc/80m5bOLFvUkDToXlVPyGLL02dY3hJd0MbCcAMkc8+56o+UzQAhGTP
k6NP0cSnV2BTUPQ33gGtzOBqaAt+7mdPmrQcK4X/xTtVNhfARMzzklPKNhc0hKDmtAk62MMs7vLO
21BUtEB/Ehdjeh60Tw/zb074L1M9EJUUs0o0c4glrSPov4PfkzcQLFvz9byZlITymX55jscT7ruR
hZF6GEaKVbkkhKCMrzx+HIut1JvUz2IRHYAREITjxSjRXvIf2dY3TJfUuhLxBQ083tQ2jtKS1X9m
eopTVhMBLo+ABTLTyIh9HwvfL4L8wW/9fs+b00QbEx4F+9dLjxAPtrkRwFbj5VAO2vGuoZSDTMWJ
oGqHFUtnSAwa1Ggqt2eedRlyxpFQ8pcbkQZSQwxKNs/9KDNlBFY+cwIMZDgzvhBR9wgr1Z6n17yM
b2hvmkjsvq5RAMcXKd7mij8O4geF8dTsUnTkGdd9tQFz4k1V9ubSikIufk4FpY76tw5m7OT7zGao
6uNkA7CSqKpgTgW3TZWdi8RyzHuh6mNjbPyWCn6rEERcjyUhadSOwHqibMStNTBQSF6eTN4PFacJ
EHSYMfgQLvLnScvZ1hEvxVcqD8bl0iXop9LBxiXaMmo09lO5+pvH6GLRjUY8/8UFMqUdW2vdMWWU
fq354mggvkqEMgpZEPyZsrM1ZmSwWyajV+ET/ZgV0YTcNxPXoEelwfwWWxEt8wBEzsva/Oeb8+RO
/DQakLld/Eyt9P77n96UJW1x+VOabMfJulKx9B1zhmLvJVtzibC2lDtG8qm1CBEvueVCk4HeT8SO
6rt8dB06xbQMPK2notvMwueBgzhbUDg2YUf+c6SuOu/gedEZhMp5DSecfW9pNvnydj3lbEE1gUg+
9jMcmf7YtbweEGByWfTmjfSPAU0gA6OARi1RTs3TgH/tzBrrGrALSjI0oYy4WmPMvNTVkEZ84Mq6
s686mhI3xehFVsX546N+45rscaup2ZuQGJ7gJ2sfGuO7GKjdfgf7w9C/qs7H4ab0+Eq2Hheb+5kl
ttRy1yJQ/Zhi2bnstc/s5lqn5lFBbtPxm0ggWX+FQ61knMNh+2CYGvZrQd7EuEpBwsTkwFspMX/B
h4jzOtmXhzHtwOteMwwxn8q1/DpbVWyCjYjLzX9lS5zu/7rxxXfSBu217ZpvrXd4UwaDIeMC1tQn
QmFTs6FILiiulRBbCUiBUMIDvghaV48jQ463PdbTVTMeqxelqc4t4Xh1lTLLcYhMTez0d+sHZoRI
mGZtxI8xeX/OP79xxlOCEKF2lqV7wefQjep74llSniP0pb48nv+ioYX6sO7ENM60w3tl40Hv3OSa
s2oq3HQX79oTgupwBMKfnlA1055PwW7GPJCgWUM7vRLYux0Q6Xps6jZNLK1VhwrYKnAwKPvQ+jD2
GUrmP8DoFNuGfjs4CW7vg2U5/UVUt4MU2tZCFjrUCrWvZ3IvKo3jXU4QgkUXxu6yWlztouA22+GS
xmGYTddcRL4JT+Jf4U8LNUZ4iBCsWROFk8siP9PWkbsrGDTI6vX9X3hD7NwWKe2f/mn00Vpq2JAy
Wy4vjBmD2CWvQbcZ4vPAHc/WD5fvxTZC61zV2y9/HCKtmr1lI4LbwhpjF2FkYuwpSYl+I6sH1UYf
GoKldRAVLgCRArr1YZiTgh0MbjgUdJPRnF9LUsB72bEKZiKcRAS/OucQIV/+j7UYHhDbNl6pedeD
+fR4JDQsRdP7f5jgD+0rxZ18UdB3p4jmZGJ2tn3H43qoKfNinO2coUQliNhO+7jV7goO5zhuP6F6
+WtyDKroCrhr5bcWYaJLFb4p8IaSc2dkBxTlRR+Sp2NdYJCFWAqFLLGIi2hhkJPObNS9RujuN4x4
yC204/qfgCxRbeW8A078uZYFruTdGyuVFTPwPR+zxHiDENSciBZMT13NXSpMSTzl1mcMZvfudb4j
tjD1vRnUdO8dANaCfLZeHhsxwZqYfVALdFS0HkK57fNT1AMaga8G7nOtnGP9v8glj8F1vfLGaD+y
j28ddnr2g3uKqdkLWjIl0qT2P3wIqeZbZdeVLkdRKP1zNz+3SrwAbkcVeoqSNGEar+1GJg5DKYit
hj2kc3Mc6ddDOe2KwZp0LJMbkHRJnnhbGg7nGrIMdZtBd179f0BP/ZGyasO8z5Qd2Ey16/OECAoU
zshDURyb4u4EZgmkbai8EQu52+JLW58o/hl0B8Esp6/B/ELno3W6MuyoD9zmoJrJ3aVg6GvKpRdL
KabJgRT8A8jwR9ZOR2j68cS7Kwk2eC0XZDJ1oimvymANiJrz1yUwynjG3JKdKskiGjPr3VpUy9WY
xHCMXWU+TD+inhsD4MFG/x7CzBUWmnKfE98fOj7m7nkBUkZWEJ8ZnQ8nGZJq+n40jkDYEfoqp2D/
FZFxKHCdUsVemsmY7NuU/oS0L2uY48apRldp34FN15ilHUPQyKwVesYTapLu0F1048nFoIrq9dUV
k2op1nky7ssGJING8qaQQk3Yv3lXAnmihrh1+92CDE0pjX9rKhvjlbbtYZz+wcrCe/wn32qFwhpH
hzzf7UdzIQwWLRQF+wnnFXQJGbKX+iy0KiQ7rd/EyZYjPe/QTKlnX8KGK5m6eDE0cKhLUFUqyQmc
MePX9hLA1AliGo2sV+gDuZ+GZCInGf/AAKfvQ+dCdiLXCy4U7xKDnSoXNEkjmwdEiH1Za0rZlti9
Y27yKws3Xc9FTOaD6r+zyAAH1CYnc4mzLqnsZAz98tE4YqDmlW6YA7hwif3Q6sXj15MACrByDK/H
a12P77p/oiuOzMVupW0PHTkQFsmjbXM4HCml9qqVaLZSudfgLTGAem6lsXTL8c3QjpqIzZN+8Eiu
UBHCJUQ4pynOSyZ7WDW8fMVd/6AP5xvUVTLADrCwHAyRBN9COBSikrzAK7frt/GMenC+Mes7+uj+
/zhxpl/KE/vCSkMu3pby67Ajxm/aPYr1nUGeuttZIm9H77xIG1xnQl8xgZ3xvXXZm/j9gs401tqL
NzBSiwykD1hT9YUaVgttUqFjVJs+cNGtrqYMdbkBKMRDqWbLlNH+owhYq15ao9RFCDE9a1MBAYCa
u2LEANr1ACoToxLBsNqLZdi/eGo6dsBtkhbYW1RxDfU04u7uTc9Zpufvk4VV4PjjecdCU9CRs+ns
ygWmbWl8DkQeau96Eq84GDQnrJUxs34u5+vrIdIOiKar9c7izBr9WsKDw8KpNWXyZNOI9sRH7rxl
MASL6m3d36/Oo0KR4Uzg1OYPI+WtWUU/pdEZHaiUIcJH8qKidp1AyFvf/x57V0nv+aKwVq2byn4o
oWdxoFP7UGqaZAK8lUjjhZCuubZdixvWdwGwLZNxMKRclpTTkeHw5GVTKx+FPGq7/tjelNijju32
aP7JKjrZOhD6npUInCMmA3hJrou+SThsScH3EcrRyS/O7su3nEviCJNoxrrOSf6vzICnNGVfbpx9
YVx65Dd6nEHUkPeiG50/pm2EqSSq8TmGAQGcUyaBehYiLcX60vs7nGZNAPepJs1iit3zj8d6+PpC
HKo2mfX26lng3zZfjmf6YbGghDzd+9ndprBnhSpfAuovMGjF6RfjCDa0wbEvNvLXw83H8wilue+d
AXyNlSFvqFEbLTrDPhBp0iILzbHt5CqfojrjmQsX4od/Um+OT7UxGP6hYQhWHAO0ynkhVVBdcHkB
zYCbn7Bjst41WnrWVsX8PcM1+wVpCTAZQ5+LczdK1+bk0j2CmNAdRDqzvnVxRiNhvSQBLm4/xdXc
4QGj2s9TsdBq3U/kHwf4u3tbbm/Bapzc6b+7XQ0AdGn7T1P90dUrApQq31UO/KjVKs7APQuqsm+k
ZPTCt1w2ej/nXwPsnaGxBa5FWy/2LkeFNpU9FbBmyeYh1Y7pEVVn7FV8cJIzjc85Sv80wdv/zOfh
NsPIPPDQQOU+J7l0Kc7yFKv+DDOTFKdtYEboOgduy275aZ4/cvUQD4qX8JxBbPup8LX8U7OshVGK
yGjpUr4bTgRjVK5JTv3Gv34WTo4kWFlm2UNQAXpNuTNFDpHqdFHIcJtZe3jqnv7YYHD7KNFvJj5x
o7n35g8eXRQBeTS1lfMIC4iSAti7UYyODPDNdNg+KJDvu7nwJsWaytPEqXRgjyIyuYKwSgGz6Ipc
hqejzP7IuhX8ow/GfVj+pJFxsQjssr984FbChzMEIrhEi2Vaf9DliBRseP6oyp01IqOyyM9LoepT
acmETsEULFzb52vlUzsCMIsEQ1IX6DJc4m6n7f7ttD3WP/vBHKym/wkoDcBkKm+3xdCL+a3i9+Zk
KstD93tJEXqozoqgwXwl5B0i90XdhBoKS0ZvQdQTq/WM0glo24nY9H3lHnFR7xNV3GgRvT37H2Eq
P1NS+2sMjfc5mxouTGyE7TTN8VXZMGT9cBN4jdecAZEhZx1Be86hIND8+EUmcUYyA63F3k0NLpmA
4qpGZIr3kVOivMP06yUYWBiM4g0dCLQdsqTaQTKIWHmyiYOsPOLzXB+PzGYvtDL4f7pMBn3uX8zh
2vO+Rt7nvrx7Tz5rZ621P78dHe5rjyKKG0yZ0L8zR7Bb59cqytJBDNIFBoD6fcuywukBYdyeyako
2pvRTE5GbMEAJCXXbAjYJXO9kLt9FkS/viP4WGm6jIx5QrSncwgEs4cIZBGw3Mmu5qxO4d2lrlj1
fC53IymRP752V2rU69g21ltjYNMe7ohqg6AHQqPjetb5IJDBQ36CjlWNqJdI5FNdTfbPOq0jgtvM
LxxADJGHZBEXK7y6a3/gYLQw0EylnMP/GZIjpSr2e+2ySxBIRTXBgjxKZuLQB3dr33LTbCFR9ZcS
jorQjwKSvw07RSzGIyv+/bmtNQUXvrqkM9kB0PDqmbuTpXmL6cdFy6fS/XjjEEiDdUvA5A2KIMNn
PqkL3TEgAfmj4KLKGc0w9wMWi2ZfzMgXec9HjbZRgHlwh/XSCA85dQryy5xN/UZydBXdyDuHsiIz
9zGzeljQi5rcYj1miarlk46IE9a7cyNcZcQG5k0ZaoyYe38xLyl84smr7pG2LnVbRs1YAwHIDgR5
sVUYoEZKlSZXnP+luPHi5AcT6H31n/fx2V9iAhnOLqCbb/SibRFk1LBxFU9YiYpdNxxuq91nI9Wx
P9d2rphNJlOHAFDnJ3t6sjo+Pdv/paAupn8wldAT0lVz/dHYgqejX13Cl6X/jRIeU0S/SZykB2VW
nhTW6CxJFMrCwLDUexvJ7mZodoWlKABaTtZYCm9QlwB3lWnXmeyfWIRsEgK1uXiNqKUCnPtk3FyD
24ri6FSCpNkaD6hUhJknvpR2/yDOk/iKJuLMXuPj8Q5VpwNVc/rqMbLc/QdXpaVCWIE2dBodF2Vg
w6rE1GMZspu//eYC/p594+azlPl6I0OR04O7Uy+BB7Mf5Q+WbrY8n3cta8mWvIVAM/LTEGCqT7Gv
lP5zex057RilV9tMSQHaF4DEw0Ykv8832lWg2GrhKPeysrKZLQHY7yw0xIc1eLHfkjL7s9VLyMKM
CIB8HHwnlvxl+1bhCjwmLcvLlNrGTLno+yqIwE5Y7q6tZ2jwmgGwJswG0c0cDZc3EnqHPxF67N1o
8XKCeP2smSXgxEFUiZSBHZPpK3JLiKR7gOp/vKHVgeyUvB7skaEG9hLFfEzeOzYQz7rzQHD5OtqY
PHxwO8K8edB76UxGib2zUO7tz8W8/+jVSdyJJZuXtpMMIRUOiqJufusJWC3Si0sIUoDy/TTWgQ0V
W6+LNMP5cQuxmel9jWC/0XZB9GA6ChKkqywvwq5KxocebGTcaymmrkVTmu9i1t76HiSsJ2HVCMp+
q9Wab8d3SLjrKygeQRSW+h8YHNs3m/voCdYGUGz9PMmdA+6LSf0jylqsepRSEDdboAkT5xrWARC5
FESIcp8rBbNjFY8INO8Rrw78nG8pDe4EO9dr31R8tzpB+V1LFJ8PIE1IzHJbg96lb9JU9TSi4w6U
BzJa7NU/D57Ug0zauG3Vsv/Ll1pavhZGjMNIbiNQx84ucdoIExgAQ2d7KGZmEzuAyaEZMZ62B7iY
mj2Zw4PnNIBLQUMYh+z9fpt6qpN2lTve/5H+5kn4/nJBzNdXaCuhLgmxUDCOMqZ0QwfvbXBMW0SN
EGOjPLak7go4aygEOyahrS249H6G/DfWLUvnz5Y6aaw6PaT7n3qMOCLXPIKvzSZ5567upZpFozFR
X1I0Gt7auNt5UhxpC16J6ozE9ZfAnGadj6bEHYTC9naCn4+ZSChK95WSw3kpDPLUSgu6Zf744vhs
9tc9v9ugiHIBrJNzRF+/IFPReA1NoNDMTAU4xgg9f4pDNnL5fEhhFSqu2KwFXPz5mlAgaCaYNVxj
afSnUSG0pu3z0yqA5+rK+TE7HNWb9UarNvFEunlDJHJoF5oDI1SguL16aHc7pGbDcM9E7Meoe90C
pXeclws0zfLfbj4shOL6asAtlgORVscef8MpxoMsJsB7b4SNfRSRCHqdesYz8OCCX8FUXVSNdlql
GpkESDrGzbLDbxGoEqecjkwlN1nwH16ejrzh2I2shXTEfritFJlEGcTMTsuDLSD7S3GnmANTGxTk
CyL+gNNs/DZ+AGqiqiNu3OS70rX4r281w7c4/0ngbsF4ONxZEFxt/DoElg1RylONTH0zE8eIyccV
IKwIiwUvhxTfPF5mDBY2uE8KEOe7gs2FuhDL/gZuGETDg7+UGWZJIuWNYLbqw8Eua1e5788XoTOs
fF1gEmZx/SIQ/dKJdhkon3rnYmC/6k1qf8DB8/5dFqDkaYFdmILNI4PmWZMG3FCos6B/zlAFMZ4L
MhVCkSElrY5v+30nj7rhpY/KRu/G4R4YQWN0IUnXW85aC716wsbCxv3Q/JH0aVan/JV6gP6dKSZv
tgolKQIiw/9p5Kg88u8QEaRrHsGgvxRiGmtA1A0iI2se0mPlW8N/rOFQjQGLGYt+PfKxn/stuzEg
7/wK0fASvGWPi49q/nliuP1Gexm2njmFwD77pm/Hvm4HImpWmQUzKx5vi6BoYWpNkR/JmjUdUii0
Hx491TWfV8/gKzMKbQl7ZB47lzvaKth4gasAhLoj99LjzurYQScxlhdWs7sp2uJUB5ZjlkZf+ewA
ro5kJWvq21TXZiRXM/7E3emrDCAEFcaD+8PTdqujspb4g6E9xGbSkWsIi6uAX7qiFqsS6gmReJTL
6aWw0BfeL5Yhs7qs7dXS0mAFfEdeaa5XrHEONRkG4GqqjM9k6rvCf9KdeyZhIsqBLlmHyIeXD8DU
unEIpDJIN7C/QOjb3HvdNmlEE9YFJOxmAeo78Uw8diOaNAX7lJJgtx2jkwlKUGx60k2+1cOiBnBz
7VEiYAGISbLYPQrZYzHozasvrEtgkvvXl9pIvzEvakFyziYfG236ePDwOJOYTdqx9xXDDXV/5AaP
9DV4e5xMCgKco7T6vDYziLsZ9cgARzns2jOFradx+jNnlGYPhZ375+LyuyjVhd4SnBen4OYOhhK6
Zm9gYfoUXvQyqKG5Zchftb7Vit6FykSMbvdrA+yd9x8PtflyUo1y2xNaIuAdycM3Z6rYS50KGJIW
x/Vu7KC0XhZI8IFNB5c3qUV1smpSjTgp+Gr2o+P0q0EI09pwTsSVBAmpzF7svJ6qlrHsYudywIGn
75UOg1TRxrUDoMK4KBFhHt9yrXDq61aNTLpNDAi47YBoyuIx7vJrkg3SouoZyijyf2sLB93LZN43
Iengy3pqttjjl2MGx5FuUFDZYpTn5MkKdoPk2zsgdc1FfsyQv7+2ROAelMNpCL7JZO5YkRjGzUTC
aaXwFuIS2gqlf0VVecfA+ehyWOHhzurWotoQQQlHAsY2ayPhFSjGL2nlyJqyLT/UOJ/RustyDDQX
lUo3cWfS8zdABpr+4P+rvAL1MoW8b4zZi2trHsC6sjBJdiXq0r6cayaZZzp4Yr05Tt1KrNKg/1HX
aw8X9SY1fF9PIGeX05DqwWagpsu3pQ9m92iWIrWsHUO/NU6bKAGT/0zqRpHmLe24MyT1denDe9Fb
hJ2Lb/ZS6Ii98dieRv+Dz7q4VtWamMwLZ/2ZRS+X05oLXbbRKEqLQ9E9pn7JwhRSgHa4zHH1McrQ
56VvDlsijHek4Ezu0kDvfm99hZMFXhyeYwZcpO1NcgnnfBAG9IDpHb91E3SnSTG1wnPPK3u3AExv
4uHr9+h9kHo5n8xIq4KIIm8JQj5+lED1nCtxb7+1bMoV3Tv08WgGcs9Fb1UM2NiiUni1wPcDHuB4
5nAyFNwXMB3E6lMBc7ondgKYrG791zAlIornnO8dPW37DlfKfExu8s3vBqrbB+ikp/uQvJWvfe4b
DCRgP+MFtbGZFo2EKwQVtkEQjJ+wq/+f23VlMk6+9bGgs9UfJumoEUrNiKvhnXyn835Yj8Wsbgkk
edtWlT8xrPbTZJhqtCYI8qJo4tfcu/ObmCV4VxUXmZeHfxVQ7xB2aTIP3238VBwIiTAshSRTJcDT
akGuODc5m8ln2+8HMOgK4dsZiDzctnUKSV0TWuFtb/ygL3CcvV25nJZa20AMU+C11x6GWlzyGYCa
kSSRzSUrlNwfoICeiEFQ45p3FFbAu1IaHCm8/1BlFwP1H9OU/I4H/+dBsmabS7UJfsHtFvR3Wh04
4CqWaYKMol/dLVVYXZcrzaidWdB5Uj1jZ9VVD5Ibms6n85u/ggeL8UKeiaCPTdqNv50dbt+LiIfB
nxIPR6GYfYFjUnGRxt2U2Rg2LRiV9OAbs6B1WtixlLeWQ4zjNjujk3lhSleeP+SnkBY5i3ZY3MCJ
SsltqIPsZzK3xeJjDa/37G8tybtbBSi1U7JyeiRGgPQiwpEHuYrEtpwIv45niXO7oS5/u887wOOO
x+ln8PEEYwYswSTlKM9qTXwxBiQD9HP5HTRCjNA6iWFGwOVXcpD/dQCr36jh+4M//0Bm4uG3+sQW
qS4Hleg6/jswzFZR7fbY7OgCX7WmOkvhkyi+/Z/7p2Jhof5appLqF0qZ+mYVRm/g9lJ1xW6lM4DK
lSvuTu7sKYPmOyPlECse8EcCka+up960gg5utVZMMVYL04JVYOHBMylnUuNdLLgQAlZfUToM96mC
Vbl/UQcNpnnkLto30nOrRH3DEtYj7q5Drq3JpKTGzM1mIsNhkWn0unKmSx7qa/cB16IjpfxdzT/c
lPbu8LsK9kjZO6l6GKTtXorb7jxfP717g31YtOPqni7MkTTBhiK+3g/zuh4vHGdmeTN0wHtaLD1x
vfjUPqRO50OYcZkN/5vLBxYfQeP/8Dcjix8a7GOzsRJzgLbmUdVmdBSpxZSWQGtZBfZY20Jx9EoN
k6SXsngHOcOq79d/TTHeq0hKmzPBxR2hxLO8RnyfIAwh2d1J5S1nTL9lJkmuPEn8bDVs+PSpEvIs
dAJiyZmAQ47FtH3/79rzqX0P5mkNQDgVDNGHa99dLBuLSoEwiPxgN7jerL7r+Ib7K8Fsy0qx6xRS
ZCA7UMyZBuKdKf1cZOYtwCjpz+Mm2NWPiLvATqErl7fRbHil7clTwzrhKfu0A9uQG7PSmJUE50sm
U3/Smwb5FvqfR/R2o3gNsYP40dUiRmniNOaF1wmx2iovQEOEOzVHgBBkPVrRTsCbOEvsg/VTTMIC
/LJUxI4WJVgkwjJp+381w07Kp+UtNDke6RZpQEqw6WLT2hm7KhT+89BdwrJpNIw2DP6lpHvOsHIz
yXPMcJEczIb5yFj+Q+26Lf0DsPwO5gLVKaEXC+rlXMA7WavEAtPz66fgIdzSVBZP9tBbHhoB0/Q4
uTp1+lq1dJmW9i18HFKLygGLzsDAoEw/Tw8u67fmoghSglRr3l+4r/oS31FBo9PL9Ify3H4TWdu/
d2lLj2n7yu+rSsmfZLuXLBUPsAXbgaeCHK45X1RR6vBoD5He/oYfCDdUfsXciOTFVJtGG8vturiX
QXDevya06RqoK1+MnuPhnn5jnWuy6Y4BV9FFO3xAn1JR4RHj80ewRrZICubCnBFDuS1tE8rhlp79
7/9CfgBOWKjRkVo3uUJCTFFBZjQMhJpcvzUqF5jAy2kg18ryR5I+PJ8nB0bNIq/7ncBwQkmwpfNV
EChvXycfOi47cJ4lkq7oE/2aXDBOLQ0tKcMeO2AYeYrV4inSwCr4LxIUsdk3axtWc6ZfwUAfxFET
hA4fhRxQCngzXM7uJD8ca3N+UkCYYl6FgL538msyPfO3T6asU/y77oaFy1PXCrC431B6FV7ihwwZ
N1A7tL3YXiXPatTsR/XodSRJPlKgjVK4eZWupZiKXv4yt41zOUZUwIwYZlKiqIOwpkSiYrqCDXPs
6kbVUCKU5Hj1U2QLrXi4QHUKUaInvwdRu2LgB5M8SJTpPlxcBp6yyuw0zaQlmhwsEjAdMjoxOrBA
aAX/nT8cXV2hUrjT2Ld5KPAkaMzTT9tDRl7M+O4ZdGIjq3Ad+KYIQoap6GKUjfsDXdPt31locUv8
PRbWaENCpl+EMqTMAPqGzXGOZkqA6Y6xwHS8QCT2Ce6/1Lwl+Ng3LOmTyZmwykoDMurc3WxicuzN
oba7IbOYHgOerF+2o8o02fnqhR4E/V2UqgvHwzQaipC+oxrNRg0wdDtq0H5v1XjjDmEqoniTSZJ3
10iU8qDvS9jg5CvPO+pelN8WjGrsavv2y8SlblhzvfLOifoXqhD1020FDHELG4wZEPm3Xat7V9lD
y9KifqkYT3NfIWzFUxGg2fj5DADZMh+1GqIywqIeYBpCQlJdEmfpBzE6/XluB626OHHCu4gdK+9C
y+D0y49hheRTapP9O6LTzX9mihfEG+zKzW24yIn+DS2Er5IxrO/Ui933SlIkl8GASYmtz5WQAxnC
uCwBrdfct7V2qDwURlcahqybo0AAvSXbwQqYtRwhHdgHyYAEL/un77nUrFG6q25h8N9Rw4UUk05M
eU+djMTDlzpQi79K2BrlHcqQUHWmCP3JQV5mstmCMf5d37MVvIjyTWE9CcN/+T+bBt91OyP93Diq
MT9wfKFzYSBsm821xYVH0/0Zjgdf4uy2G8JIVhKlH+tGUmWyWxPTNpZpQGTePVIPtj7E41rEJS67
WkOtgeZVRY6jOKL3TDyAHsTaL3JGqS2TjVSWPdAzmgP/RykXjupvDrJ4zUdX/jvPERc0DA3nPtZv
Aiet9dRXJrCc7uPlEDuz9PU+ms/AIvWDVBxEe4i7rXp8iejbywjbu31BjvTQbeXwNBCOhI7t3hT9
FyfDr6hbptfJ8Nf3KkW9W1+T+nO9BQOU+jOLXc5qhdYIxmPyInKYFHrvNnm2pVUQGwOmTuMHOlpt
3NxQ9DXL2gwtbtSWgFlNrWn/NKTUnNFq7G5RRhFGiZ9j9TkgOrGAIDYDOrSdAAGYp48t7ePOkMHd
rki2sJwzRoWowfk6cE6yTJGzqbRSfwXQ5vCxyppyTdRhunUzYFylew6G1dE/jjBQxKAbs5SSQ6Hv
vpGSzP8FRrAIOnX/xUkBjbyLlCupShuuJSWheKBwD0TVdFMAx2dFpuNV8kBzpVnxJm/deEp+onaN
QGvuCunpanwTFqyyxrE/oZ4mP4e7xJKH3d2ufQ4DUC3SskHOeHhlkm5APPuGmIVpi7TH+rf7RYor
Mwz7jWt6sXrBBb9zwKaGHBCy6k5N7mspxqKUgNx8J1uYVYop6P3dQ6ywf7F9Yvy5P7pDGLAqVQ9G
VC9lHT4ZhL+Kscb/aDRfL3HA2Arj8ReTcZ9HuZLRMC2kFmMqlMlABo/KKjLi+gM5JTehBQVF1QA1
ki7Q9AXAd/K9QFnfms+7X06QtBYil5hl+WtsvQucyPjE4AbboP8bkqCJrZT7BfoC95MsLtLtevv7
oR4iFjg96wi3/gqYE0K64J9x5by/XoEFeJumND2tsANtwj5cyXHeD8Fge6AB+8XrX3C5RQTU15c5
6mC9zF+2xoh4YWP8rqCKM0id8bOAcyRCQbKY7JPDUJGBgibva3QH6TL/kOxwwaYg+JSjhCb3FBhg
vut9mmssBczlelYW/vuI8sa8ycejSCSWiX7r8evg5GCpRRrK7gNputz3Z/V+grAD/swMaMdaGd3l
i1q5c4gfdJ4XoMJ2ZVAvm2lvheb6siXKkRRnaKHRhvpBQ6pYwAGgYXdUisWsVVSKQD/uaHBbkRO2
d989+begK7asbw37mfRvF2Qzx2vNhNRkXZfySTxEj/v0qDTEh2Hzjdm6zQSJ1JV1H5c24CazeVkR
SxzNjlZKNvaN6YCZGBY/kv/DA9qNHpIDT4kM3von7+sEpa+zQqaSAst+kWIbIC6DMGr4mijNyBCI
0608frZbfFic71wNTc7YVmC6XtpvttZsqnVbKbRTovrvpkb2JvQE6CatHMUUGuNr8gTCqpoqHrYX
KltfmZGT6m1qRTvPDunqm9eD8cZNDdYsRLQdN6+sexYye5v/0cftxh+MV6M9JWUv4W5b84/uT6YK
k+4hJJ6ohyFxznT3bQztgeIi5+F3A09/RxZ4Whhk5jW3ARKx6Q5ol4mk2ZbPYjX4u/1SgdvOLY/p
8WBKpILVfZxK2WPYI2C+C1Rzq/VJJX2QRLBzrFlj3aOyPglffpgc4KpHtWcq82MBq04FhDOecju1
yWjb6vocklopPjHnM8fqaeZPy62HcEKNc5rUTV2kgR9NdT3o05j2ttsTGvTqOdR5fEPpHGQEKhMP
82uGSLqIWskaUP1kmVrqG91+j0/Fs+u5gfkLbOIKDJDSQVXEzA0eRcyG46XEUlG/slHUdDH57PtX
RV+RUjWcJirHEct79GTgxotuTzx+jyRAkrQ+jxuROFZ/wIsa65d9h3Zhhea13dUhd8DBWCW/gfmK
RN7WjJxpq1Mq5bcDb9BEesAMQdirIwJ/xuqdlpu4joB7zecTQXnI7Vr39Z1xal8aEUHjFp7l6CMf
7NJ0wbo3JJJNzeLi2rYQ+TC4gznLnkcPvhFw1BXLdy0gfnySyt3usf/ZJuby+bkNaY2a1wECsNjw
Ra4ZvbH+I5WdAB/G1skEFu0fyHemZwakxioACb7yz28wbYafhe+DpFt+8jEM2r3QVWroXXt54cv+
qMVflUyV6w0mspDQHQyXEk4NisxyTpdIEXK45XVYMXmy+Q1JP0onorClx43wZQuc+uHO0LHhUF2Z
Lp14eyUmmipdF/i23dGiC4GQWku/x2fWMQqqMNAIIUQxKqAP2DdgAB3rsyVkUcP2Pyg4s6Ejrre/
+tYkipuIi1TD36h1KI+teUoPj+DCsGCf+pS5+VMTe/njIrktKsjDH/izOh0yabDhQXNwNiZcKf0s
Qq034vNYAvcegICNQAJwjxgFNGqpSF0x/GlO3qwAqMIrIugEns4y9AOgjUTjviEdX6d+8xQhwSUd
X7jj+zLmwSA/jHWxjKDxpS6lrcXLYDtpGQvBRbClOBlVzR65kfzxP0VR546CB2ir3dvkh44jS9c2
ILRQjgh638xOojFbMKUVdjePFQj+tV4bIFbqe/vY4nTV03Y/YsjD//TUGM72kqYeHd2FnHOLC84Q
nlGqywevgeZUFr+I0LoDFs68rdo9DGjaUZCb1yyRXY8w1llPfzB6d+3t12w0XmjmiH7PWBqGdUup
EU3dF6Czf4HJqSQhnUM2hQf3pwRfQALBi76wLT6khO0/H6CNcBaAwVJvYNuIuiURw80r/2AuHgtn
MsjLQPOulOMFs29AI0JOg5ikfRPzH9Qg1/nZZkMSZyJqUXS9rCx/oZN/qSQ4fkswsvMdwK9x+ioR
0NSM8EtOBKHFM3rwx/MHQ3otYc32mbueo2z4E2wjAilV7KH0EzmbhGXyaX1YwmSbGjoW8MaJeTWo
h51nuczLYiQcAey4p5XoRcur68Bu3ANoQqUal/Lc+xd3QcmDzXxF78n+RLXmbeIjNW6/HBPXYWNv
SzBRd+MYup6/2KuVD+YQQp2pBQN/2zKNLBbPf+/aWISwfhBkOrtnQqRw/rsOotJOD7er8hs7Ph4B
5lF2vSbn/ew1byrNxk9Wv9Dvk5lYZV5sfiqDsDvBmQFwtx8ftP6VbyMoxgPU9QfbhjvqEreU6nY9
Nb1Hz72RFB80k2RviKzSpmOyVbQjDSMhr36VJmjtkQk0edvJhHrzsisHebitEYUAV1/Crbhu0eRw
WKLbFoB6Cb7kr3DIi1nAMwHZgrI9hKj4NuUyzw4e8Ne6hkJIJqM3KWX1AYz4bBxEQXWlVrSfvHRx
KIJFECg3zGNRLdlUexMlgyRj6MQutEqtbEtOyvz21iVoN16IReXm3QZTWtXmGJI218HQZHd5TLiu
ziqNmyWElK+4KMRAZA5xIgwPG2v+c1UbPRQ4UVcsP8C52UnDB8yafonX8pHA4Dy5q7VpT63jY35C
0mOwjtpsIT9xy190Mdws5l30z/N3YBoPqfmaSDp4Lc8FJ/v8F9f90KzN9Dw3YqdYKp2FGTGWpeQo
YwzyiN4CQSDM2UREW8TdPgejMkVYTVPTB0etrlvCQy543AYzjSOy0w/MToxN1khX222SZvpavrX/
tVoPtPvgjFbULdWRk4U7lVdF21BUTV+gaf3uXymt9+Zr/t5iix7IU0yhUQuZkpDdv8n1tH6hH4Fs
1xu0UE2/QqXv+UD1/HH0PVtS+T2tnG7x9Cju/RBrEb5qF92mBMxuIolEJLqw8FgPGXoq5te0O3JH
4OKqT/1kSXGiCqD4ku+x5KNeIg44ZU3ekP4R1W95RfHI6cGM8wd8CT99NjnQIw6p8pfOBW0D+iWj
oVvbsdF8cqjqTaryBvRPR9jv6sYCvM0HqU2cO/2GpJyAEa0ObYgSYU+nqKTv64LkA1Lpv0Hiu22z
j/dealvWv4UI8+2x4rDiNtDBCurve9Qe98i0xgwAYLrl7JhQBmmU8aVSKK6qhlSf6QN7rt5oQwTt
j3W+DBo/EkyYFrmVgTWWLFEv7jAbQVQLwyol0IGNrCJBKkuWluAOCGFd5QxqLdwGMVjwFPlPIce9
xuvc4s+zAd9TQV3mBV6UzSnNegeZD9AiTS48+3iqWadx+ps7gzmhHSEW41qa4Ed6Tj0aLpZQ26gQ
P2e74UcrxKsfQfJdkdUz1KnL4SsYflCM/u6EaIi3Qga/K0due0jW4FBfe+IG/Dh/4cD3O19bhCIV
aX1B8bw8M39/aIswoyeDpkFFhjYClyrWPhixDLaUqjcZOi4et54cp4Fd/Q5fuX0DL/xZsRrcMDCV
yeeoifkOCylkr+4sVj6UKpHZBcRVqiDhrN2Zre7JmQ40oso0nqGJP4+BWg/fXUsKhn3JmIyjp/4N
MW8OdxxfbtWF8c63g/dnsCJbHfe9R8VdcJAh8090sKV4f4nSIMkKog2cThqfYEEfgP70/zEcxSSw
5wVp/OM0kJvwZenQ34BjNetHkJLxVMRSt7Ki+q3NzHv/yCCuJxMTD2y9uYdb56ihDwpNYc+Q+0xe
J9dS1z6cKXsgDL/biV00/AbSf72b1NLfzGz3DKc51zHLBtqdqcqOCNSgypxCFtECnDlvlCNzsUH2
W/LVPeji4+tn11IYyZLx8nTM9WvSqTlTIDwPnfP0gWhD5A4ylaGnOzCb6+wPFglGfJAkbXcECLkF
FkQwGH3EnapphZMXcr38NxhEkkoQlhj/6f3sAF647XqUneaATro5mzFAMzloe24JIZJgo5W9pYvg
wFHISKuP9kzOymfrYa48h2xSFU3avzgMIj20V5oWsYIFzMvy/WMN8xghIAz77xy5DRV6LS20fdat
Bf6fD1b3AJtgZjmhVhNQBohMF12ewMZFWYHSkVB3FWSn+v3BaAdhaA3XNbWslk04wBrb1oVG/Jn2
lB0dTEQttxttFfUpDo//53jqddpitvEcsJ8+/A5fBiyq8bTT5uRxijYLGVk8tn7yXgtOGoDVY/JV
HGHLb/w1UY6vjjU3mvgE/fJb+GwVrSXJSlMd7Yn57GL3yAurWsCB0NjuMSPkYHmsaywhPYLElLYb
0e7sv4Us8tcwvaRg6LQcM6IdbVUxfeCU5F3T8CHIsKQSZ9zjxARDO2f4nv7dsQkRJbeOGjHVQ8Sq
LoMfJpLMtJX1E1/PIg8hur46z+WAlHZt5jK+Q+AnMZ6s1kKpy9ur5/0QYaUM6zD7Kpw7VnfRvIk8
Q2keVkUcGBxw9P4na9baQumH+wKh2ZKVIlNc7LqHVZCzxea8cvxyNxeh0EYimCLsUA3HQzztW9wk
0ZGACHM1gYZg+q8gcXAnkoaKXuQtFr6ZZ4DpPTJ6R+4Fn0YvcDttZsHVeYDikTVKUJMOc2sn8mw+
ExlkLvOz/hcOjNzHjsFK2ObRjSJ8Fdt0pqADzJyk2MZ7TtpmRo9lAz2VWVm7FbGlejQEcLStC7Aq
p06ouVtYqR8B3bFzyXZRAfqeR1YeJqNd3asO3QXQMOVLe7c0G47jZvkcQBMu9dY+Oa7kOsHqR/KC
q2xpJuq+F8OlA+1bfi5K3PQXrGceTFgYCsStoWjNuQWKx8M1KMR0R4omZToSlwWqddGSur8+N+i2
vrnLDRSD+82K6iucyyP2oaYVFZYBc2NemuU1BoJQISfXh6yhmDDgIKPvltA+pyve2RyHnNfVajXh
UflY7vOOTd434YwcjTodaBwCsyt9UmT2erHGWD1wWpJ9yOr4cEdDUUkCew9UppXP6GeNtIy/d96M
8/ta4fC3yetgVnVMmsAOZsO3mHU0VE5zswiFH9nVsccbT1LHFlBNuMr2y9iVkEbDpG3vq/Y324Yw
hV4sit0fzJCnYjzS7oL+nnZ1pOa63Ik3U1MYZJmTZjnUrh/oUWKleWltDQn9myiS1a4kUa0bijM+
wz5H+K2uAs/laM9ixsHJ64MDyscbs6n+rFIIGaKbls/nB9mLFmCQWz39Z0V8YX1ZmpgfP4u1SC7t
Ja3ktzBU/+bZ32rytCD7O+BR291svp13uStQab7vrVbmUTX7AX/k/R6bI1KnRdWKoPnTiZb2K/nB
DVzLEX6+UitWLnyYU0Ys9BZeukOUxejN/xpozPh+58aSa71Dnz44qZzhFsu4v/JZDCBuryf8aZFH
CGBzq5gkxIGphNPDzvd6sokG9kTDzGCYlmyW2TY5aKX+7FZTgJM5fr/wGNB6Uzsl1jCiljKo/zxH
xZfDD/sc3UQtX2fAXUipS07BaAmU7qNYWLZO3u6lupn3rSl0DwzZFKVsND5cfTwOaYXQbesafLg3
AJD3Jr5d3EAOJyTHuBfnDiHFC9IQg5zULW1arYGZywAEmZ2m84ru9JtVVrGIj5Z9V76Lz9pjdONq
sa6jSbbiJ4iGNzTxuWk3Ha5I/9sAs/YKJVrSHjcVuoihPLOK3LRP5QA07GEZnKz4xy3jCZjYwnh2
YK39CR0n3llJEOZLXOc6g8Z32uXkgMRYSqtA0ohkUdV0jfXTDKBg0h3ziswUXfhjICUvNkD9iRhm
QbrouHxhrkCuzIGjQZW3n31+kDWzCL80OhrffSSTjLjIRqqhOEy1rjWZbGE7OOh7v0KF7FjubThc
KTkUZFNeO1kS0r2XFilP4LU9CHVip6Kr3dyqqIiVeBMl0TeTvRzvqY+I9HuL6ypgzsAdph1Bfgkt
tpCgkwmI9RNASgTGK2+kzWcbEfzuRvZyNgfOC9wDmzfPg4eOt3YJSKQgxCQ/Izn2U0arO7DzD974
zlQ24JH3hEwR+8bGfYPRZAPWJIOf+pyWehTfNNkb76SPfYxFg/uYneuuBf2KU30s/YKVn5/g+5Hy
kZwjmFFNZUCo93l+Cyo5HyJS4Jg3aSm4m25lRwYRTMf/MaJC0j5BwG4UKbNSAizDpOhFAb67Dgzj
N85k0P8UVPX9E6Ax/EMsxppTD2fIA57RIo9rmv4QDYUamvd9mYyIAx1AOzcYXYVeA+9gkJiUdc99
ituxlKkoErpGbF/mIvAbw1UQo6dHO20wHNJX+qHWI06c0C6AIb6dQSDuh9Yhinv9fU6DjetuODMT
rwqPOw5D+skhoPv8va6eGlw+zbAfsVR9j2j65MZeqV5gTYKow3zoOrcMdJtcu52nqMM94C2eM9iP
52Rwy0xMwZpll4KdCNTyFQTB/Fo9iCHsfWpHS/JTqLawA8OL7ZOGMCwUvXzxu697Sr23qCv3YWvX
bO7H/2vqvIxIqS+FpVIwdgpixa8WvTebTXV20/LH0WuUuFOMkOfAjs3xtVl0g4OlVslTaJ9lh+0b
Qdrq0G22eVBG/JHEUefXsDpK1t56LCLiLAPV89Jp7JoDFQ8iruHH2qWm4yD7bTRIfJ1dxsP0G4zQ
RkaKVeaJK78cmFwo3x2hzPShi51yzwK4RaM/buaemejOZo1jT4gnWQrXFi3Hke+VISEjJwAgyqOz
WH/Qnd8aqAdCR6o+wF5Oj7Jo4gRC8MJhtASBh5xDAR78suA84HQQGRz+e3KifCVwsyYn1+4i7iUV
mm9Kq6Vq472lE+ebVuhJhjAoh8epEcX4kjqZOtlca1Q8ODLtRaQC4kC2/MxYZxZ2YTbwa52wVmny
l9ZyaUPssBnxVB0h6UaoFhWcbQvj/WNZcHVPGfj0DuC8yTfhaeiVaz44w982jWatw6ivzXInued1
rp9WCk0d+71dfT3AzIdC1rFqx2qRs5F5VkviWvvW5zgqqCkms/Bd150h6nMKj8rHyUiDkMZyMIgW
ALq0MY1aCqbVIrpRV8o8+ROc48KVFv9CQFe22V/DK8AfzAIgmnzxjVUtGMn7KKo2HgOkxLGEDCyN
a9cYP5PrdyMyLQ5SfrTmIWip64w8bQB74b99YMRr8fdcQ820NQtQFjWRFdJqajuZ7V7wN2kJE08U
nYAVFzY8tassxMLEzUWQXJ5Qd9714IcBi4YfIkCxRFIdAtQwLADuP/7kiV9LPSwWKFqxEeYxTefJ
WTCMI0c+kFauo8aVDYXKXnap2a+WozwgRytUYLlR2L1eIO4IVcoPXOjB6Ue4gPEYIebXhlRCHA6s
sHi3YJcgJBI59+wUuUe/nPEWdV0uvoB1hlcVrVU1SW8ZfjX0G3z434oOum/2AtPmZS2HmVH9EjgI
MoRki5t/2ysFJwAQM0t0iRpQlf/KciFBRnWKVOVnZvA6gOw+CVH82AzbEWRg35Njy/Jbb7/AzMlX
rsAQ5r3wEKPHx7U3VAza7TDl9lQepuOwv9CD3yp3NvB0SiZ2nzW17jZI7QC8yzcT/rdcrCoSr82h
cHgxXIu1Cy+XWC4OozbDZUt3rKg4WmmynaqMmQloUGdROz5FLt7ta9B61ugjXkJif9xAj7fROP3d
A7AWPTNKFHdAK5n0L1svUlCkp9g0oGZ/vWBwCqERsUUx0fx2jeXFZdVRmNTeqPlB74K+TtSvfIuO
Ts/txbsewSrQzR3xm7PgHQACk1kRXbSv8JIXXLtGW3nyT5bj6eS6zV+kkH+pVpmRhaGDg20R5xrc
gVnk7Wp2lkIrQwzaG4PfrArtKTuR74JIhJjVnLDr84dKA0hL8sVx3qMEikDHrTs6lvSSbYZPZhtS
uaCja3kU41IAh2f4JcDN5rXs3yXGggSfvYrp/n+0CiFu3FPiuZ/xXeoM/Ul8x+Q36G7t/us1iR1z
outb8nFVtW1LN2su9tregyuaFTLsW0qGl/Mdp4pCVYoyc5LvL6SYaPoG/3QKgU/pBW2EKHlE2sOl
J6GLzba2kssg3Aotnibsun3XiEYoZxkOJCctn0D9Q7ylZRYiErx7yU99YAPo437KVhcwiF0A2dBW
I3Era3hhb1SfFnRlr3laWP4Q8S/yeljFDD9x69Mg/xJnQktabR2lKRVHBEd+cu3YeZt8jeQw/l9w
/hUplf8wvZrQkoNuShSUiLpM9R0Hgik7bwvX+7YvyMsgiLVmnY7QuRlZU56X34jdU0oxRtpi08Os
w5EvBrbcKgAwWjeBzOQOZ+1/40VvcSwCEIozxJKybjfY1OBTdaf2X9S5HGyPdVYDmKAvIf+Y0odc
N5/VPjcQPfaIIgOvYiZD3+2oayWOnj5vGya/3zyxsGOojE647FusjomSMhqGg4z3ZdR8m1Rf4cZI
zE1BQTYn8pOlq7ffqVdTgPD4DTdqK8HtfYfj/Ezd8RdH2tiZxAvqfM9d5gKLRsXX+rxXnTW65QQT
WmNUr5jvYyFbH0WDob8r4E/vuV4RkNG2f3HKgAyjRKXHE3r4eUJHwoRITA/R5yFh3kHaYocSIIdE
yirhTybHTa3nKqwb27aMAtj7N5sCDTTFM91lkl27kmrggbKERBx0S07KNIe3zNf4CGRI6EKGkMom
XkI8QbRMDO/foodX/MvIFWi6JCHOaA5I/80/5UZT8SKDQg09DwEhtyMwBS8Wiu0W8Reb+73yiPUX
xLcDZkKUCsewqhVcYX9bLc1pOsokqVoWxjAAqKSEf3W+KUo+cBRqV+JtphoKGDQirCihEX2HmQIg
NWKx60ZodyuzJo9ZWfUDLabODY6660smUnQqKswbXF8pa01TaHXe/+/CAr3X+UN5z0CC6iIdb48f
QSlUgKlOWuk/pkzNWYB8mhAKM5Xah2p4YoaRM6ZyYClf1lNO9nJzisN7GJ7P/YDRlXM2miu3IyY2
AIK9daz2yWwPjHxOrfSbeIXY3PT0h9ngWB+leuJJjYWuACeawKtPs+kuQRT6MtkcepeZNQ2YI0It
yznekpD7E9Zxf1QkrfE42Fcrf0bs9IWn57ixvIOl3dYSxBzxrH2iFJB5dhGOi1ZKIxnULV6c47zz
X1dwDgg17W0y+SGdIlAEnjtrFWG2UiqhNiijcj1qcTs8hdNJ8TLSuaFm9RkzDDsGVltiS7W/JsiS
zrly40mzeD1yLToyZqHIgutQqCii5rAgForVeFyPNKfVPtC8HH1PpwIMfT/IRqof5Dg+nzfvzULn
Il8fzu8jkalQVNLv4f24oCo1RHmWDUt2Wjy5bI/gbJ35iYjJ/p6DWstWdOOADqwDjFZuk6Y6xha0
qIw7SGifZFGwH8tqD06G6SwiidcZ4qNt9d41S4BIDrkH9DMIeM71TU1+e0dZVo3QZ2YxY3nuuZxb
Edq8SjdrNAL0u0plHRgrHGQoOrdnLAsuQvsP7hzFyxSnvRqrBhgZHyi+PfzQ9hXjb95awq+R+MoY
r6po3xoindZRMxu/tyYb8GX1vJWh9Qk92qFhTiE8JjiGDS19maPV5OoESDAkr0a8H7EW6X29/nDR
OzuSxdp++bfEUVHJV++LqijVM+8QHL91QD+7AxdRYPUL7hIEZdAxewcXagj7TZ3l9mZmsZ29rErY
e7c8aWfQNnLSpRPXKDYegLUaRMYqQGhSTzh12r/PArqKg/zdERUTHqmQjYF5dKVo5+KzKHR0d5L4
MECD0BIbQvNGF3fWo+aVoO+VxIJ7iLMpmDJULunPDcCZPOisITkyoT5XKwMKgrYNM2erW4xCbR72
bRhktnYbwVWv5qUZABzKZoLwhCM5Un+vvErgwHzGELT6up71FI8G35flgcttG3qsFyL5zxqkAmhg
F7Ft9UF3vHMWUfZ+Y6LcBveIuiQYtYIIdumJaU4kFyLYvEDbr0Fq6137m9KDUy91fXVIsQWY6xV3
SdkDtHqduIoaO/fKIn42sv7rnboUna76qDxmGVEnyNuWkoaavfheqoHSJfjpwlL5Sekva6wPuEdV
0sjPZ6Esc9sdIW75gS4f7YTWyX/Ju7sduLRy9tYkqbS6+YHqBMUTHnBZRHTXcwtpWTmyGVcJC9OP
kJvv2hyVTeXCuadkJFB90WBk6lDBl7oxfNE2g+1bvwryNsYTTjt+ksao462Lra69tcKYzhkn2ok+
LQDRA6fJK/4YeXHQ3PGacf5WKlBmXf/4uMbxW6xkf2ODcO2s9WU7q3fwa00wQRqifR4ZoxTy6pDp
A2BnHPXEQDzD3RMZqdgqA654NcRmy9WWkOPL5SnOMr2KblwsXja9YmGfFllzFEAOKmEkuDs0XIWF
tDtqDhvcRr3vTcfNcMXBlG63qz4qmpMF1Huopba6HASVCZXxwiZtsyB+Jk2DGIs6VoqO/hQrpYCl
xpxi5P2X59akqYmcESnOtSZdXHPci40F4y5Pfcn/XSuTe/vFLoYZKvxOwssl2vN8cbIwv774tLoD
ZGtBulS3/QUKLjV6uRwByyZR253MASA/OZd0vvpylJEaDEJl0IUhwGpP/GBLCWXPPDn5QKgS+Q0X
cix1c8E/pNsHy2GBw3TtUnKWO37JiTNk5vx38IMaLQmbCk6cxx7eMJT50WeDNBKLPYdCivfyWRR1
wPpMzv32y0Q3Dm46oDedPXIGR1c2WDLYrSeFAGpTDbLBWQONRDTGf9QVSDG5htSu0t7PAu8qRbud
kyDhKGIuAwaPHgcJiiwNkF5aYP9K1Za/av3OCFPbu0qEpvHR8EIX6Ia6EqeScyokwzeywVvlZ0n7
hM2X8MFnwrfIH54Tj3y9aFkF91BJI1y5vLErSdsP67ynzCQaokznglib4vB3ybkJ34VPTvQSMspL
LAkGRaCVYX2J8vNR4j0HPdMXZfNK7Y2UAsu6CiEmGnRHucpB74PN96HrKMRzB6pxNuwPDMQoXYEU
AQh6ky3Mb0qLAx04QR/0AnWhJEt5STxpCc2haG40G+OHa7NTRoT0uAo3UPIuuG9wbD2dpuzWOY8C
FA5gYfE2WbuJcIRwMdEirTFmDIdY/dx2Bi9O+hfPN38Rz3pWlyJfj3S4CqKFStZJyoNq7/ajFzcv
MEW9FvWdvwvKnJ6apBLJXd2DqBxcVd9gMj7hbsWQSvT2z/g0librFh36krPNWPVbR1sH6F/7r7Wb
NmWKjqYGlv38rJkvBx0+Uj+1NRn5iotudAHihpcjA5bNd9+mvN21RKkLVue5Jp8s81agiuzU99i2
kX5vW1eJ4iQg0Q+HRA4VlCosJ8NHzWEL6UNPQRtBMZailHt5oT6cbOArp+m/Bnxcl46ee0NJrvTc
KoZYFNmAuIeFKeqA+g3GVgC3x3QNcxwKdQNDYxIOiiRhF4/1oAHlN1TZGz+CsNun+XZD5xnYfZEp
Lc+8ZAFYwhgeGk9fsaEbc/cq1I3O2GaB6oqQBOrCU6BEc6F8CFX1HVBsCoZZaq7LF2+pFQMB2OG6
zXEdaXUHQ7yWDD7C9AuJJa6wq4SibD9wLVUHjGu6vABpZREB+IKLnPV7xygAldrVkNFeniXlG8Yh
EN6cR08QIDfFVqU3xFP01EmTZ0zdW/3naaGcEHvVLueGQjUEfAsiKDEkw75KT0WUAvRUrymUexnx
sFi4bZ0gL10+9ETDU1lOo2sG8u9tsgTo9ETL3ARSCOa7OeZhVbp+bqhLKpcCiJaYhILdqpod69dK
LQwiKo/FZj0aV+5GrLS6U/B8AzbpW1JyI2zVW5SZ2la/oO4F5jcqUhL03YAfiHMwtYCkWukodU0g
FpPx+7GiQAE4v927CgnEsXpIlJPgcGZXlPQV/zIfrDMBCvo3GtOisfPCdatqJQk1X1Q7psV2SJOv
wk9vi22Sx2TuKYkCotARRM0Eu4ABgw5zKfarDFnXWVGvULMb8a7v1EhgpKVapSpCnysHOFKKGvOS
9P0VYIxOQCHgPpmiAuoD2Mlhh6K9nbD1dmWRsq31BWgYEkP30l92v40BItuOKxY+Pe6Ygp01zFuc
w84LZeLIk84YN03Abbdn7B2ts5gho6YFYSIjDsEFlZVexB1xgoKsRHjemGWslT76lQ6LPbpqKV7t
97xBuuve5ok9l2qEC5v48Z+EjeLLPVzINnThP/EZXwHkQ1y+DBvAaEh+yG6ghhL1u86S7/Rw/J6+
YUBZreOH/rEUJvOlU8orpSLy8LH9eWSiswsrLaYcc705V4NdIn5Eqo9HeFNzE6fDdTwM8NZqNU+d
MCIu5McnOWESXU0rwxLcwE7YhHF5et3f+RFehZIuLoTXXeBjEdRczgllcNDK3LthYYq9NLumVuOu
KRMBuj6Q22Fe9a8hNvJ7XAKaAshOBH6xaUjLRdmEGZSQMJaBRdR0md8xXDwq1klXqqK8p+CdGlWB
lpQTWAUAXVJdUqssBETdhAsuWmuXX2DHH4NYApP0YjGa9SUNmmGrJcjEDgjsXN9vxmUw/u1AiSJJ
8FxItykPdJbtQVPBtZKXdAf2W4vbsQoCP9+n+dI7fbsKO547tFgpqKIFkkPi5kAHQTNKlTVLGQ/A
CdflU89uQQdEZowAR23Hef87OwalHVJFMRIwedtJMht3ni2kgbu0G+gB1LgAZLokYws17mKUxGZt
SROe3coqUh9Nbl51FwZ8VLsh2iNtJ/DUxUQkElGUr5dbBjSG8x+wmJNjyBZHML9ILkOrQ7b1ELu3
+reqldvkPb3YKHQdcmnMq/b+buUDXxLIkvzLvxw6qLeBXObzUDDxv0c88lXtxOXxMYTtRbPRpHEg
Co0/n7t/BRsGKIiwmhoxWiqyGZh8n/seuNIjVcxE1DIP4W9yLp51jAcA0EwoliF0tnrZeWrMClE8
jPi6NTLKA6SaPAhSITT3yGJeoi5rL5VSN1/vN/dV8BvTqvDyBZ+U+EHDtsJRgV1fjclFigLJwYLh
uI/ENw3Eo5HT12adOjfDys6adnVIujhZBTFCp3KeZB7GnOf6Sa/uJLZnKMGIeqTvlUd8tRxbirKT
WI6l1cvsJfrXdi0K1+Edg5FNnkR7qJPZAbiCVtKd9L/Bml5I98n7EnTsIOwGm5Kay4lGMNXPRpWp
s4z1FmIfZP9QdRqpUc3aZx3CIWmw+lrjnO845k1kDTeGGAEEGSrHTrn7c0J2g0qh1d/6aFcJAd69
GbZSYMIQHn2RNy9LQqa3+OrHPB4VjjG9lqXnmEWpRBw8hM0IH6/mar9kae66NgYxGwIaoMFT4YpB
DGrD194FpIm70hhMO2hF9puGRGYu58TI/vdDoGdYT5/MEcCv6bLWgPSwEk1sLaYFzye017NWrRGc
mEnR9AmDaijNJdbbwJE+8GDsZNA5PPrvY3XOWCsHECa+BqrXH2jiyQgommez0NAK12SCkK7D1LNH
d9MNEkAT1LMCVEZtDvr6ZZzvb/pT1VNKAIe14IFn4zSRFBv3bax8V6QWQpncM5FN/baCHbyyiIgz
RttacAsJGPNkLja3WQ/6OawXPTKZ0tjsg9UI73dJeMD3SlrkqOSQm3gVONvoW4BhjbsV2gLcMP6X
Ft2R4d1g2t0rOZ4/h5Xqzg9uKDqbZ6X3bJesWrBgO5FP1SDTo4YRA39nH9GfkByGSqQr1aKKHUdv
mT/FNdWA3IZlHQhnMsXCrqdmkmNifmCEUWDkRs34mgU30xxrvGpwLOfkcPri2Y2qBmMmyCqTbdoL
T9yV0bWJZdnQeuBHftcw4lGu0DY5RCBdKgDQtl9twjWSxauP8OVGwEJC0d5PpuP5FYvX+nanRKMh
Ourkdzu2Znlcla7hKFXJlnnaeI879MokapjWuVM951n0cqnjrG6RifjlvO3050VNg/+V2VxelG87
1M35hjO9xAf8h/FGYR2bRG6brYZWJwU7rkIZTnMj671QYHjFhmn11BSGhVLAScmbltUybkAqKcHw
6vuEAGEXEbaw+Yk5vMcamhRxrETpx3ElFlaS/DwCAXNE3eq23AHHyRZUEWZUJXkH7XVoL97xfNEi
DzLL7ye0km4lujtqbntvGGdHvcZNCw7/nZfmofARCZwlnZ7WMFnswfTzyM3toO/qkhARncJdkced
tukapbiRWpa2AEqkxGqlWATHUNZn33GXY4MKRRf0APsMLsoJq5ify0CIpcrygiZZ7a59jLXXWWZV
v6hP658TjXwysLSROU2yu2T59450ETBBDGPdFDKkzW8tRcPLILfh/osWaGWpg2ipEyza76yAzDTF
LlPWvlUyhBtjShrqS21KllM3q1onWgGElHR5pbx2XOI8iyTj8k0DDuNEwO/O5XRtXrHUrpplM/w7
tbASMN0YNJ2XfPCGlLCc1UkkyF7kvHmbaoTw4Hau1HF3s97DBFYzP/B7ZASNKYSWhW0R6neSLMeL
3JhMBXDnb7vmFDcSjDLbyf5nSPR+v/BFoB+JKuPMIb965z9QqYUv27tFPN/HJ+EajtIOkZO1XQkE
gjsIIaj7dgbBwe3MuHqzJKTQCdxCIJIQ9aTs9218P7g3/UT0cuBpPOAVE4wkxumMZwH+p3xcpXda
s2xIaQCA4dDESsWE3Fb14p2gsSVvdS01ngk9ETkMfPxcth2z313PG3F9/g2EgUc35ZZpEnAyXO0E
21rMjr/sXdCGfHHMpl+NSuErsuwA9j1bZmRyGISllH+2SO1wYipWEYJCuweCkbc/KgXtGHLwBTfE
DnKEcN2hens799hkTq5DGa/VoUbnL41Sy0Ku1o+3JCpITdsKkwfHWI5n8MhhZ6YQxHwOo47dfper
P+qrFX9dijr3TNznuY6foaWGEAsHN+v+tlMHmPuLQtzzoLBFxn0LMwgWSoolD5nlnw5trJHHp588
trnzb/K7AuC9O2wAzHDxddchNUreHH6R0YhcZED751sB/XlkAgF71Cqk3mtNJpJTKlfVZ6O/0YZY
tvzQ/u5HoWplQ4BHW4i6KQx/VW1OZfYUxqmAJEeybJWJGvdFKq7/7UblBUi3z3zON65u2EYaCLgJ
Qw75I33ls5soFPSvgXJNAjywfXGu8X1BAYw6aUlNcRmmlVV9+XEsd2v3h/SwisIfL3uG2iVckwna
rJwDgruuu6ALUipFo6+oG89CZFiBfTFX9Eyo4TXDBF5ojvbIF/PWz6m8weUVEP13Uthl6NmXIvC0
/aiwyZukkBEU/JRM57ULRPSgTPzdBauzyGZslRpCX3wTCVlsRkAKMTHKLgzaI5tY9D9JPYx0HcKE
Mbh425VbIcMJtg0RmAhv/+iV6lTOhfmVDGJdEspChaJvV2fRsDw2reacCH2yJjvShJ0c1PugZY1M
nPcET5L3fYqAQJQxFasT1mzEHs/MnsWZ9hmRu3ldzrJgph2hSYmI68IsHY3HdQ9QcR0oJjU/2C5P
1CJWW05JcRJYEYseHMlX+S47blWnuJoxgcp/GSWYFR9xitznuhG7eJG3DRSWENIiZgoiQg7S9SXe
AGkUDYciKCHb6YouwwteoSFVFPmMcXPlOG1Zqf28imrpMWOnIOjyxekaRJZGTTPCjRoD9QtlbYS3
zTPtmodR1gi4pPNWr9+6ZuQsVwx3lRC1MH3X+nrAZq08oqY5QIik+MfRLpTksRsKQ77mCb9ZL2Rx
BcMJWzisy+oAcl6RsZEsmo3BC85McRm8FZnOeWj9yBCE/uVZP/aONG6q7vIfcsJ32yM6+ASZdqEE
s+IJPFKttLqkvP64hJiZff7NHQdC6mx/hP8F6dgbENJcvDoNvbDXGI4bEJn6ihiuVHUvo1M/3dVM
z9S6jBWi6SC4DJcHLsDZ5kVJJVgs7lIb10fwQjJRJkBoWGRO+4KZqje27g8KpEt4+8iPo4xY7FlA
UxstUCP9PKuDYiftX9ddj2ty4ESINqgLrvXSFXu3h2lG9dRrxoQ1ZsH79bl6QN5CbICaHhR5LJ/S
0LXmZnZrKpoyeQ/WHKpeH0gTcjVlP8XlbKTwrmiWABu9U/mNEjtKhZM1Lkrj1cKzUerFj5hfXnkj
R/lPMyzMGPDWsNpY4iWilcMshs+4BIAZ7IbrhB3BsKK4IuxWvMKqa1aNkHCWo1Z5KLWuFvQSfltR
xF0d7QUHDDSNIw5KD5alXtGSTcFUVA1FEHMDzcXC+hgG94RIswx+W5XCCu9Cbh+NhGe58e4HqsuP
Jnrm0vmbhfv4/DrY0Iypw4i4gPA5o1r1tMS66gcSLG/3hSf/4XLlyzVFcgFZhVECXX1OInG1iSg8
wQvhaA7bZnef2pYFqnFJs7sA1nBbSd/9RHnlKLQ9Gxt4hxZ4Jpt3WYaUjfd1Q55tEFIdZRCs4wiz
yk+gMGr/OoOYFFfk75O6uQRNorh/s4XqFAivyoDpJKeo9ubR+WjmBrFTm8NT4JKFVWqFz1euHC/l
83LPbXwZyJA7+S8WNOs3X8PBp/tirYIHUgHZMcbbCLRl5aArLJrshMG9Wx1YZB1r/IzdGZQ11T1N
b4wt/zn/F3LMsxHYrWxhsGhiL/ZTp+FN21chkyDKGgGH8SpScVu+HALN5OZr488tSHVKIlogblzg
YHX0s2JPMOEgUnZzuG3NbotwCrA+f5IOvjZgw5XGjBAXYEjD/yNFvyOBqQlg2Ykv38avii9hJLxI
Ra6niWYE86zJxYZJ3DBR5kruszvohSZ4aIjwW/r7isGtDiPdVqOCr1oMW5o+1e4bhboYoJZs+lo0
BlD6aKrMAjXnyIPdoMZ/LcqafxMC6kqdBxYvd7/tEteulsvfgsmY/6B2NQ6o7BkoQR/qU0ivlP5p
9ldf10cx1MwG/eRDCRi3ByYrJCX+AOEp60tm2FyED8b8FyRc7/0HIJtLaPRtg4QTXcjOoLWWKhut
QoE+1PvgZJ/dMB2M0l+9ybbct/fyYkxZRfP60xNpaVb/1jALlztKoWMHE5m5GReyf3Is0uvHjZo2
ATpDBhjIAx9ne/L3Dt2tRc9FvcLswo0+b9x0UEtQQ8Rp9YJRpeAePuJyTcZRjbKChVCWlvA7oXVT
uDOSyVXzBwk8MvzFTrDJUfigQg7OpADeQoz1uPyKdbMU/eXyZ8ZYDaxOSTcGMULoNfO5rBy6FYCq
Vtx+4IcZryT/n6kRXsUn3gEAgnx/v70Waq7kkxBnxLx/4kRUHDr5NAK52yYkFBhrr6c4tg+ct/Q6
wUY7IyLFlwWyEdehteHOgYMp4XzYep1C348ANDPApBAhc93gJkeLcVt+MQVtjnfr8bAKe5FljKGL
WCMSXZUIqEyhomDiwDWbf6xF/zJVuhzy3p/vO+x0RmvffVOp7bhpoytiQdjVT7Q2jbGgelicfIuk
1Uy1hZSoQIQsZriXY9rgMcz2BqG9wFeGPJuDHPitndVP72p/smREZZlb+dfk+zNdZDPe4JgVfIED
1GKP4Q5rnqwaV8Zo3wQSCB56+i+orMIErcdEcb/KkRi9D2BTa7OLpX8EgH05AMavPQ/Dyuitt+wQ
nxSclBoOhEK8b5f5ffqRNjKuUImGXiR/knMU0uPft7MFO66rPHXPx8JH7XHYNWhmk3PL33YRiSl2
0voVkzWebBWpm/F2Fq7G+nmd92Knpn4e27UnhG+kQfdIr+CDxxoC2hB9nL0PfqT5IZjdh2NtlRrO
cysTe+mRGes7lpxxFc0rUx6GCGbS97QENIBu0LWERoRhj8jVHBweVPYjDBOVmuD5c1irSXZG6y4G
DA9ToJ1jvYnNp3QsLVU6sX96MNq+Gw2lWy3BmWLEL9hWcmDmGVg9H+AzuU+xR9XJFOCmVnXHrE2E
N3vp2KN8tEjBDCx2NKxfo3ro21f5nF7SAbkZHB2cYRuTfKvQVA0ZXLOOMEYU8PStUAKX/rnoYD59
jNfSmrbp3skO4b7neUcq96aQ/Mxj5aWBu/96CtuRPANY94L33uI95OyY1QL+SOaJANGregLa7olZ
uVeFhPdLn5TBzwbe5WdQ/OJ0SlTVH5jVES5fLAOIijTAjjc/23LD+KNeC6996uqoddnVUpHBQEdG
Qyol+8B0eG04OGbQxP/hAALDRRhXezdNIqd3z1B2Tkbjfl28Vq2Pencf94NXqAvHFGvRq89J10Mx
bBLlDov5EfBb46VJeMNAh0NhejFOdRsEdd1Vra6+abPo4M0rTglqF435gFoxLjd+rEltrKyGAZVz
2TayzgfKR2k75NIEfMt4pqJWVtIno4JHHHJpN5eTlPqYjT2Z3+KShM7hv3ULZNT/4mjEgoWxUYK5
Orfac28JTDtlMYBWSSt8Nx4Y0M9Frk8zsZbTghz05q+TmufD8P8GJh7LdWMt2ud3HDn3gKYyroks
nU0dZoVkD9zGjOkMfaaZi5eVP3YerSXvhtOdvDiIYv7eAoU26WipFHciqckYxdM8/ZnPVVQJDjs0
WyvxXJqYAAuo5mczzR/CV9ePc0QfH4NN3Bp2VKHSdKtdKEotEiYFdiuFH5tcQivqp7jMFTj+5qLW
pVXMME0OeJIcCheaDVEdn2BwQsFIOTnbDeXeVWeNlCmS1vCldhR8FTi24wOGlRP7V1sfy0yDW0DD
Gt2DdI3J2ZEyUx7Zxq7npSGDwOCasqomO/ravGWp34X5CRaASvUqJk9C21xryk0SJsnPF1mvPTB1
E1YMaLYJKE4DdfvOvwWqVkKzam7jzN+vptTji7ZUSaveXqsWjM7UZboXsCxKhSr0NE1UIPPPBNgc
1PD3g5/uF3gA6ajefxXyB4gnmnCC9sNB2GOl89E+pVFjjbX4ocVWh12g4ASESxC9e2Op5nJeONnj
7GCHl6hVIvpXuFpzQrVwK4wGwhVMHQKyrWtdeZMcy7hO5+LCfacwi6koGNh5cac2N/j7Z7RBcHXp
PpzcEGLW7VzjwNzgD4J5C3uOjb2QEQKi3cVh1+gOzPbLKebNYikOmxFBQ3sODdcZuZfaax1RrlJh
roAnYfxg73dwDw6dzOuBpGS+dpcpnfrbPw6NWMwx5dtni7yWhBBAz7QBh3MoOFD56cgHNgeZQ2bw
BKPUvbfiZPaslzgJO5vwNlX9zA937omIL7t4c4225M5ZEZWtXsWg3WbrFsTYf3n1kRGfGg86o8DN
J+JnZpVqHqBioiT8BjPuMzn+sVfJmR2chgcyvvOIqtsZKyWf6jcNjXGuW3yeqJeBgZjC15OEte4k
DNVVHzsGswvc425VVNGO7mawIPGCsJsuJOcwwGnDNh8oQL6Texg7yl1s4p5VStpGqXFN+sBX2YWb
iGNDW0X1G8X7NoreB6Hg0Tn/PKUNQc+Ssi2Musa0CctFjRdVfzZeN8R+QEZdzWZu4Q+Ld/TuD8eR
fLeJV9U/sW4Gm2HF0o9mtieU1jxYdz/54zD1Q54c6Th/SOFKPjCEQP1noaMFB7shpYN+6Oo+RBV2
/IL6hRzwYWFGepDbxN689Re9nt7uY2lJpfsgr54ILvLdDMYmMzE5CUxErtskIZMkFmpWhgRuXPBU
XmUMtePJC7yUxYL1DBse3NzS/oKJEsYYIhwCH3kQNAOjldWwTl+U/6M2AMw9D52mmbAG7CPdWjm+
wLOjsF9oRsReYZ84zaRLzolUM9Fju+ba0V+oHnbntsVUMxEG7KsfEUIarrEDRzB0ZBC5rWwploBC
y3NPgK+/ru9H5Yav4cSSxFzQKgNZJ19uCsYqwlG4r9mkvGxzDmH7EB3nSc6jFlslciQsxvLpOU1I
RavdZicJj1KxH0OFMSO5MUyBYeyTc3Oodqr2YK/nQdL0EkkC33+JRNTRfTDK4blRiIdWK9NBTI6W
+WZBPawQy2bXl9ZMLb8e3Um0/YUQjzJvwK9ZlzdVDCUpUOPbkK9Lm4aRXHmjawovC7FLypgJXk65
ZfU/+U0yn6DjFyllQ+ON/E2NziQ6b/zYbPBW8dRzXm8GFpYzfushORrowJ4jlHOEZfy/kHzBMxjV
uHkuz2kzL7qPYPS+bgV/NtYeA6acG0ESoVdsSCUMc2CsoddbgQG7IbGWZOc7jz1v5DiqIP0ynS92
wxyO5ZUQU0tqIMrPn1ivLC1qWVb32mb27LYLQlPYl3V10AfXtnPrvmva7WLmY4MHkG34ayNhDkrF
GruSSObOVK2T0hkrGZDbuGc3q+Kn5LqPCD0FR+N1IEHDpBCWrEAyluQjcRDfTBs3IB+eZEWz66Qn
On/Lk4Qk53XVq/GLdofuhPMbd22IoilHMKgoAK7FWSVxbUsETAqz7ZImrJ/GdpUmSa2jLkF+g17T
buIGbERVwlUFJrlhbkovMkpZISYDZHXzTWHJLSZDRFvLXhk3eJPf9WccfwFFV1VBEMSjR3JErBa7
vJLyAkGeyEO5Y64B2PjXx1vQLGzBeG7+9Gy7ir/BlLIew7yzR1uZP9ExHQywCFNFuJftQj7MV7Zo
KTwznfa0FOKcETpWYv4M9FdRi63flW2+e15oHNjWmuzaYqzHtQdLmUwBHinbJIKCJxnVviZJ978N
KhBCIPtg6emhraIp/fTZtiwXVUQT1tRAx+WtH/drJ1p5fXxJ9J9QYORZi7mCwsvfWLH3l90+uT4k
TiOVXJrbZycoiOBG5GyYNjySmjiCFL5dUfmigzisdBWe6E/dnoK+X0tgc9u6m0zKlm+p8w1F66wM
Ir8T1aRXyjjBnNoSvRkmzMemZILs4QzW/C/8fEtXntxABQ+uIgp8m6mM0aH7AQFGWcvp0MXVh0+A
fEuwg4BaANgP/jAmcQuHCAHEf6vszvQt5WRPw63lqg13vK1seslYeIGpvnsVwKZ/8DydvTci26xB
xdWIpx8dZuwjMNUu0mV+LJMKO6+zvfoPA8l2O0gfzSMCmsgigYx9UVdKKCkkZULrvmAXLTJtLuYK
byAiIdGBG2STtGZ8o/0I4pCHPdykGCZfJg1mJb76VfuwM0oGISbahEKYYB4lMGL4zZX65Btbwa0y
8aJoVaIJz2G9ecjQ9VG3ug37PbEFo+J5trd8cx+sDMpcaUecFELbPODNzBj6Qr2h0OniRYlteP6W
VB279tfiBCMGgCvgcBRyIYBBJhQyB9WqXDTo7nM/Q8eAAoKqJSLFZpuhc01mbXuGhVnJ4WfSuyP5
pXaBjrcr9kVXTnOXSKWmmSJIpUTn6ITOc+ERNo1hg98wTCUG8sc1rmXu1EbfM4l1f5ebnmkh1Vm5
p6f2GpM+TNfKGwZF4XH6YF4D0BkOQqHsgwMKTElZPNecUBEKNAP48M0z3aGZgU0cC4G/DGhzyUYZ
1IM9JxmU2kwx25AgckUaPBSOmPrADPru3UWrgaPJvjTMLlgeeJlQE8LM+ZrEhzK2ikEDGGhxkDmS
E70esbB0jtcggZrI0B+EoA/MaOH0FDGXZatOOeKiF/05MaOc6dNkG38tfwfER90w1nDgetW6RVsW
Hu0TY2419BEOGXZaZDEE94Z/+P33mYrPzo7d7PZa2Z6L8en31/800y/7eFVy0HCAmZuGPu4AEZwR
tV3KxuAOsQMqx9qFZh8vpgdCEmTSEvUtWekrBEPcYM0cUk0gAY+/mzJe1PDIhAfa3F5rHZLIYjTd
cMxtKyDM8t6ic2SdT3ZOOMovVl4dNtel9sdu+cPiBhOM9iG8CS3QO2+YfqIb6uHMnp5g8/CnWjWv
NXSVAH963afm/BeyFi7oo9BrnoBxOHy9XfzdTjS0WSUd95PGJz9t8q6XT0q1VVds00vU4Tqutola
YqTyIRAMc1C7Ys3m51SLgRZ2zsx0v4eyThU4yw9vjoDzfH+hnfKjjCz4/ZTtuTxHpZCPs/VCkb5S
fbn2b+RkArkEriHOy/IZXldXn+s8i2KjavXyjqPOXoKP5w7hWHy3PZFJ/+KkolxS05+DZ+qnpYDC
n8yF1KVR+H3rI7lKuimaD2depzweDI1Fbs5fhu9pz1nrfg4Cc1MDJdCcGnkHtnIlLV+gf2+PgdQu
YXPLn+7wXhs0ZKNKmjpxbU/qsvd0cyuqTeaby69P1H673ppAXX/rZszoNHMrJDV/khqqOQA8xFiS
A9vENlckgoRuAoGsuGORKrDFrJydZf/GTkJwBC0xKhNaNiaJBLTdeJcHs6jNoPkJqER8Vn4PVSaS
ZyzxrGdGWVjLW4qqKOJcGxAJjUCUcJns8s879eYVtTXj2IZ2yFeMgcYqIY3rfRyOV9XwV4Rv5mhv
BbySerqp9xMKAS2R8VNLxPD29cncJFhU1kItMIm6F9KjBJQwzX89pJIE83CwsmWMpsvgLzkkGXgZ
PPlQle5AkDqz9dYGKJFSZGW+oxr+c5yNt+qrCJrvLEO06sZeFdwRTwPOMkfR8nM7h+rCCo5lydB3
mFJrrwXCBQ+zZGf9AfSOrhuUhrgcAEyRTLs4cql9EoMRC7zch51AzW6TNHRJYkszQNl2yBj1rjbY
F/P3uHUzG6LHwbQT6+D0HI64xbkNuqichGaZMa3+kzlXBm3MC3X5dADKkr+5bqLHn1Gmt4qHH0IK
YTziWYWAdRzgocgVPNcS4AoRw2j+elM3GvBQTfEXEUixGLXchF1tKihpTVlgiz468PqRFziC+LCf
Fw9Gkq7UMZathbb37YBHnfUqSeN1mpjkX5kM+CBBeA4LkdzrOoBM78d7YMUQSFlGhB+qfUlexwIC
7bDgIOlb8kIx+3q1KM5w5G97F63PF0+MCJTdfJAZtn55QipTqPeGuQdg2tBkNW0+sU0Prig3ySEJ
GpQZbiIeUeZErDHFyD8TEyrPtzOfWHTyHBIxqqGde2jUm0w/Ip7RuORrCARr6+7ZGBkKdh8junX3
pzGD6XTpNJZNaspzmJI/BE9SYIYIIsLFg4q1Qij0q+EKY3zdFLytK9rpzhElB0tiGQixZnuVc60K
36JgjkmtTpz/kriPb8xzzjhaTSX7zPVPKc/Wvt6HS7sVBkImWwE4PmBgk9AezAASpydSGpqbNxfS
5wZYX/YJEKyz+quE77zC7wuFhuW9zq9ZmfBSt+xSIyq8psC17CY+iB7h7GOgRTu9Bp5owZDJciW4
BIrKmNmOvEDh6PmzIzPcmhyS38pL3dw6/rb13LcyPVd9irPqSNQhNHAJExZ8Nxm6H1JBgp4TB44F
r4+5pjxkK4L1wfEMzA02GwgqUd+4GdyRtpxDoDtUTVvKQr/iD19VckbyLX2NfKjFOtHnH0HRR3Eu
MmRospFjYWhSOvkIPaMmLhg3yUYURBWKF59V6hyOdtveJ8YiZx+rAC4D1UeMnusBEVnAslKlT552
RCnxWDrEnFgUPn5c8HuRiVJoHrubBjl2VLQ474I2PTsaSZLiDL3tueNGIlq/WwBotA8Z4KJXkUad
b8VmPWcxDfB+HvcWhi28GwqsyfJ36RCFF4XQ+ftL2Mxthn3pDrwx7ITcl3oD91ZCq7aBLYteJ4oR
w/aJ37vh/URFuI1ZDTcD/JjHIXXT4ViHhbe/FJhZjmUwcOJ5LVLwqkfkyUlOR1lhCDy6bbmMZAJe
DryCuRt2/S+gkwNWUcTTaCnMjYLXprUqt5gAcSPlGd+tq7OcoKS9sxT0G8loERPOK5Vw3Fr4f5oG
dEMhs5Wjlq/VTq7FxgXkEokaz2obeFbOsNvGyocqc3BBPQk2bACWOe+o29XzYhNV+QbKB59vG74+
G6JpW7YI89ugHfz0YstkGH3SvTe4QLCiTTftBTc6Fc/zvuFqq5osF7hn+3JjLIva8PVp7eh464oM
d5/Hegj1X7cNar4uHnMvXGFLIqpdvXoxiAFPrVblHHhbHYi6h90ffxyXwooiWdYJbYkUUf4peFJ8
dsG1CjGt+qJePCeEXE/uRvayu6cx7V7bB3ZOFL4cuqRJnQ2GCs3QFYX9jklAsmTwt5mp4ESiNB/M
SpDhJEh+nSSFKc10sXmGwSKl231+P1JbfEBd7SxCDLpF0RyZSyk3Pp5FNmw24iVrLkVL/I0CqoAP
rWdzqEBBBOiZmc8wE1Fdv7pSEf7awUzb6vfIofmUkZMHbU4YRkYF0kIBINFlfbbNXP9aKz/sZA+P
EPxjiYKDCD07Yt7koq8xF8B0QC7rua5NvPTD4NFZq1FVGUbwNqJ6h042UIqk6gyfMM1tBNMNq2cJ
SdjGu5xJMB8OBHpjRQAHxiUR+IySC+WtVpQKwbKVY8IzI7FFNxID1vwmW3E1FujzFcnvAwSlma8b
jJvc2qYsWB7D8BMM7DWstDK7mX3AfGEPDXy6epGsHv5Sr99Ej5WW7kS75quMfOGPYtX0ZaXLZRs6
+DM63qh3kyVTBgJE5oXvvNKW8RXFgp5gkMT8Bfz5FnRG7HYWpTN9F/Lo7t8jAap1EWzt+nowMoNj
aLoaIdOaR+aK42dfHGMElVShWB+hzPcuWwCU4qpRo80nAdWl6rYSK5XF4WC8SF6SIAGbWpZu96Lt
IKvcaxCCQwq8blGu/kdzOSeFTaRJCK+Mk0dtJLPUkJ2QQaVl2z+VfKA0bwRvJ4AwstQqSaLju/0F
9w1oK6lOZiKmgFRNVp4huKu8cFlr+RhLwoj/phErtoJTASuEaEMNMdW/ejGFLP7KgwtQjp35F15v
GXn65mu+HrphELBUWNhYURoctMEz0eufANqP67hnmtfcS0o0f0tE1lrI9KuCScJHAXKyDfbSg/w0
RdSA86+wt1fOT6yZfmBt0BC8nDZ9NoeU2fWTZaXm2sGUJyu6EaWe5C8QsQZ//kGdMW7F3DZaYBhO
sey43OosUrx9HvfIARxojQp1SMEig5jqQNWl6nX3UPo7WIQGpvQRn4ahDhSMDC5M6z3iKgPbUH81
w+kmnx3PKJiyRZZjkkCBnRHHku3OpaHkBEgtwWW/XUmxldX6Ezmalw0mriXU5Y7ukv0AhRsuK3fl
GbVV9RWHeMf047+o3IvD4jYVSwHyMLI/WwA9nuVt/tzPjH1sQVhhXObqznbhYz2fe/CGDFUG8g/5
D6QJYaCYicKP8jwb52QhOdTwEZ37EI5ekIDw9KsSWn7foZOVJ0KWidfzAJTpyNKZmCaOma3DSg7V
cXRiPKTD4ppek3CuQrFsU1Z4GGrfgGI2gwcvTnDSLjvH5KA4L8EcG0xNMqRwErorzuwWN0dd/AN2
e2cuJUU6ZflGW6AuUH0sRq76C+0XYo6alz5qJ2FQKyJOFQJht9DEEzfCO2Vq8moWPp4V0f3QveDf
XgoU8wVyRetppdunJZBOxeUzO7NhiCLq3Y7r7ltfV/2F/3LwkNFA5Y0rGlZZZOrNc9XTeMsus++D
txO7yl0RsQqGYp8W/4vr4f/d+BWWQj6+Puzqit20kZHC5YrGGjZ7ZMefBJXCXMHF7lOqhazQV8fp
PDvWvE4aa7Sla7GM9xSj8kd+wzsMtPWnCvPjInQrgLepgLw0vp6DhCAEthqjV3aWsUYDE4CM2ueV
5RdRQwUHBtVBnrNfLq3J3eoIlawJK4IJNpyEz1obQi2ctJdXdWD8U/mjybXpIhqDV3hk2i8V/5KB
SjH6a07FIxY6JQRQnZVhgwaB7/4N71xipLAw0nrTCI/ctfBKojM8K1RvN/eMU+/1rTMPhLJQHxqj
gq+vLmoV7NJovKShWQE/dWxjrFACwgECCdo60qiCPDWIzoygO2I8xAOU4BSTVOxfw6gx6zb3XgTs
D6HKw80m6PgoSZ16VrcLFqPpv7sgchZo4ePkxn55wLhskd46dZXKGIwSuzyMmbOC2LEtb2CxBuN2
/X0Hw4D9QhF/YoAw9wIQ/inlYcaSobP0Dt2ouHyIuByF7DLJvXbRBcCyB/XGQIiPeP4WLEoYAyBs
Q1x0+ct92FXkJVBpDKR1vf/03pDEoo+PEHRcnzDP0uhCOK4PZAAbC6Fn/Iq+cGb8+EmIxjdH+BzX
Jfoj3duP8oCcBM60wdEJJhONzlkTMYKh+nXPK6QoeH/wyXqf/T4QGaVElxtWLJBhVp8LQwcBMTu2
7zG28vSl25yqfR4/Ic53B+JCc6lEDKE4+3UU6IqL8ksKOslmIuMCyOwmkXO1HcZBCjNWgW4Qf4/n
kdN/SHOlnTwQRUBcneGBKZVFwdALtloV5FNP7rreqgh5FXH0V33SCMyrz4EmFoM12Qix+9A5obyd
Thj2CaSjgxCumaCKhYptr2pIRdoczMWCmYf9l3FU0v71NchccWaPqMhjkP5CPRAJMvLCKI/cOUOt
/VL0FHoiN96jhirEXjEGYhph6ewzWbCcK23mi2VHuNCE/GZe3ptBuginK1gIRyMGSOgt5+5WjRUA
N9+lTBi1GyM9fK5DvI4ccT4rPvNCFfFuTyWaceQ8kn2NxxQnUDDfPBzlPTtkFlLEnU7AeissJxXZ
91xkeQc58tUhu6VWkyzky2SxlXBEKVUfIeBX7KfPQReyLEaxu0b/16+Oew1W/WqipV9x99iih06P
qUaJGEe4lgLUitx5AOZQR5efZMXR69PXby3iUNN5XJQLi0CG/hRKJH45s/gbZh+sRo3SozFe1VI5
xuYGfuMIsa35iMaS33WXihAyAQoVOCImpwx+meVZWrJisRcvvmVpZ9KB2tZhrLaR/IWPV9OqwsBZ
oNKri4lGOuz34K7ROXj531GR1BG+Ykn3/D9v7zV9H6LRj34p4xIWRqVmnc/6f3Wc2pH/tE9zhMeE
uL14STTExag+HapV5nU+mACTLPKolokUKrAGpMtWG1lG/kQHKInUl3fTtS9zJ9XS31IByQOOykMj
EIzJq2F0FJ5KG6p2jsIG2i5Ali8DY6VSmTs6BA29PVicXquMWtPeBCehheonmOPx7NR+Zm2148hE
CX9gH2GsM21DLBGoG8iq2TF5maHF3i7fQ8z2Br4syTzkHCOM5coFVhdMRCrpSS32i0Xm6+6Ql0qh
WrGL/5byUm13v/uAApbpNXwS2POBlb2BkNhBwEAckrIE3MnSVOVMVicRPphpr0IV7YLV/crHDLH/
ISHbMLFm9LswXCLWm4zBYKpIiFxYhn/ym1s6jpjv82Ct7Xs9kSd/V7u1T/EMPApI1hgNoHkbyZaZ
aWIm2cB3lU25Jd4pfNr3T0otd64OlrfwIAMYeNZHI86OMhpQrp6QqKNRw/p+B2X3p16Zp3/yehXG
I7aqclTbr1UYDMUQCeA1LVLqTosX6bRvbTxnrtiM1JnDmozQcWgUZ4kboIim21xur5h9JU/GmQMh
HM6L5fDKFfTydv6+a6DsSaGy1CPE6tTlHDyGYaVfR6xCojUyyo6EJEhHxoePFwvO48PnX3NOPAa9
Mb37nSa9mHTnSoTo44yT+6ss35dwTnD2YiFOZfZxDmwngLI9Y67ObnZ5z9ctnMp5tdUOfowI7TMe
so+i8srbHgUcTtwcnC4f7rmxYIZRzSARu5kFmKyPZCVosJozVEV3DgPogVaaNWI6AZzUmlvUsfzc
I92vsxUKdBbOPc276C1JxLJygGjoIDg+uPDm5W9l9yxIlN//1agvwg309jLaS3iptOcyx5moo1cR
FKUq6F5IQkcRJQZaPMmmXk6DxbCghtlUY3uCwmlCoRZmxo408D2TgEKW3hXkybVq8+XVTAyqDlZA
j/HZ6FaFFBJH8I+gpIIilvG3wx3raNfgUQl5Zm2hw+lbV5N+Auc3tpoggsgPNuIJ79PG4saRUX2o
o3z0NNDsyCeXPSQhj6VhFF0frCG0ikygj5xZOAnEu/uacOsQsi+ts91C/1NSytYa+aqkszxKnWWp
axeqUJr6/rCLCzTZ5NOSOen3Ov0PXwAJhu2ZJ/vDLMP5pNN/P7WKZGbOsYhMl04NW2y69J1n5OOE
+dcpQiWwuLHmIQgaCYDyAE6RP18P4wuWtUCVcDgzutU+T7if/T1OhCv/aPhf86hWz/Gs1kCCnHNU
rnqMYBIQGxqtLG7AD8OX2Ao+GUVRDHWxzdJ+Bosrs+4f1rv3BEtO4XeIYUVefWtaxmdfGxAlqGb0
9Jqlp2g4vhBkApnhWgFofapX6wwRS2nALpaVYS4e6c+8eNYQOJ3h1gsUKIBydV8/v9WdYu4Umo+h
pRwwZXaSg1tRViKEVub1XCIIVGvONC4k8WQoL8Bp4+z0CummgsnQFbNzjvQTD431+Sh99UW+UgeX
imZdGEQDkb3rkAbbrtN7Em4P9h0owhMA/a9rf/p57LU3hh+xITxlrEUr1g175xM8shYo2gWXtptL
n+bQPShAIhszVN9AsIVmlL1c40wcII6xVthV1QUEYAPNZwrXpCJ6DlJj+pNJoyH2t1vbtsbXsX86
qUvCqDNvoFZETQHa2PFSY9aphQ4msXWIjQaqU2lz/NEkHsA0uBAsmwx9HgotVWxxF6JKy7VDxBRI
2Mqynogn6vIMFB87l07mcnFliT2c59tm0y/PhgkVO86RaKScozQfUEth896N6KUcYPCBfVDGu0h0
naJ4Y1VgT375RPY8hT99mYtipxBw5hUMnHQSsPWaLMF02ZXB1/44OH0QdxuzvSjUVZicrHQbbdh4
oyt5zvAbp+HXRPC505r3Dw9gc5ugMP7x2axoMQ2T4COMCoP6c+ypEUzh6ucL9/n7GI/G3WIk/laK
XDYs+sfv+BYLBA0UoNkiTOcu3ALn4HQD5WSFfU1XZVSaTdcOygnBEPORqX+gf5ir3FutrmpqPpP8
JT6FBu3HQbd0/oDHxMstPJaLg5BtQ/ImmaM4SlnoQSyeq2oid00FbX/Jm6njXBH2dzaDhulEaFiO
mMg/+kyzjF8gPKo4msk+ZogAVE0AiJnhwkCjd8YoFtrWXRjlOxh2Kos7QbDreykAkS6rPyCNtl7n
n9pdGWyaGR5Xim3ZwxLiaTyLTjXrTZIUcIQ9bANApzp08lasUQ8J8JHoXSaR6XGfNKaY/tkXwXjI
knW3nPmJXnMB4q1xGZ95tUDi6yMP5BHWTxxs+3/y8uh1HSLGzSrcX0ax4FLx6PXlHsw/dnxRlR/u
nVEXxAvnufyCI6OrhOPAWqYddWEwYrvsSRgurrxTlW/yZxcoXz2xYAh9K4sfER8cOmTRTKCG4TAG
R8CJzwx9GNQIuXqKreq8fMhlTDRFeybKxPCEN3PxJF758uvB6RHVxIA4JsICUS6itMYKgtgWeViw
YHgJthTocjyflGdPEsgnnX2Cd6bkMJlNtHBCUoUlYY2OoGqoYNTZvScklI4nEU6TrPuV0m07bcbI
7iMKpT5S2t8rkXb4Ty1XtZucO9imIQR0TqgV2ARFK2k5YF7z8gQjDUsQgYB02hK8DAXc2XM1QDp0
qEQPzER5Mu/Y7hVDS6g2UwS3YhM1CX3JGvlDLtKLM2OgO3RH8pNdJBwgsXykBXqZIBqXgdmdJn1D
nc7f/dNfAoERoOWKKqmIsKUUCspHcOBpgBlYjLYHpp6S+GpnGcvaBWlAXfL2uLIxbJIzu65jnVzv
SATD9jvoHOONZxOpyb4hsP7pjCn32TzZJLyJhtx+0Dtp45xqGhKt++dmIyBXJeXdZ7qEb1ZgMk93
tf7caWbZ2qd39bXmuj8R/ggbMcgOEm+uxWcxKYtcGKWJxPqGe4fbm6xbW8vBGkYKIudP13C6tOcs
/iD6rzlUddiJbhjX/n7MhBkhfRq/4jmFZ5BcPS7LfHhj7mq+TCsvzSHVNg3JfINPRz0YaVSTZaYy
dkFgdULEJBIuiridXZjpL7GkAhm+OCNGCjLUGh0cpPaAEvK5mglvwMrmMCvY9zbJx3ExSVPLobPc
KgQAIjGtOiuRvQHBaFzo9GqsPlHsrjPvYDjv0Ykoknw25uTnyf30cqh3nrYjUemhVrOAa3+OrcX/
SC1jNFa2JaPHoo0OYOIPP66CM2kUsIaSnfSR2lECAJjsGrOy3xa2rTX1cwQpJocs/SNuNks6a5J1
2FT1ePVl9pPlk1P19CbC3EOAeqpiL1vmIhSArN1OM4qA86kefto6COvVQUDoNmszDNzcNdZoLE6o
xnZNCvahwxYIgGfBPrNtl8f4yIyDqIGS48JbNPpxbMEzSHA85Moe6ewCFgo5AK5tu4wEoCF+Bn/F
l/NPQ1obTV46jgRkGxLnfHaOOXvFzrNnELzMyAhg9lfhD6e8TaW0qXNeRNBGYNRKa9plaNUJKTcW
Tr+4NFStM0F/CooFYBVLMAKnirmlIOAP3QLNPFYfWotHmWExPpK1OymAT27Rc913KpAzIrXrykQ7
33H1iTrGasxPBBIeaunCTUxag2rSIBeYeZeWrJDH8uUNqzIqX5qJexnGTnDLrdCsgfTzMMD4CzlH
kPqhUhDkDuYWn+PtXTDJ7LR5QWmEFhP6FVpaVM5fM1X6bovkleNZSPCiVpTFa52ZGjBbAjyiOSNG
uno7vUEtyFX5+TnoWvT43ICjnIE9sTjhsBsyGYeERhQ6pIDEWQDCT68Yf7BvNB5e6ScslHe0QxXh
6YBjoQQa+1yLzWXN98BWFcYqy56/3OcUTNZJ0nPA/n867crypZu1L4ndkIfW8UvPkHfRpRw+3l4q
5KBqXH9Vpo2fFHRYxeQiMDZ3reoCT2RvnAcu1HWWL5c2eIY0kRTJZZ/svTcvtZJNvVmrNnL9hpFd
8kr87pKfCSr67iOFCu03rT1Nln7hHjSxzTWgabKX51d7WApLEf+fNWXKOOt3+Si05q7Yeo2PFvIX
VHzZL0nwAhPPBFkvh1GClq4t+WMwBuYCDEpD/N3Jr49yWjnK5qIXLqJNNXRUWXCWwFXug9yVYKys
BBgLOUwFGaccZqWHpSnGaAn+lyzkEqsFZelmdqzfhfv+hwddi7kUYHGTNADf4fBnksL7WY7Ho8Ee
A0c5pYVCfiRdrOhTEysd0HJInoXUlC3pUU7NJA8oG5NADsidyiLg7vo4HT2Ou2eCuf++JnY77gDM
wAahiY4D4u0x64Gkp4P4Y4WZ+DdJgxAgbq4e0wcXdF1RisLgq1tj12GYfpm2zMwNlW3nGyZ1yNDU
mk2887rJXuB1Ctsl6GNPn83U7BElClJUJ19rhXUXGgPno9jgdnu8HTAQOChBE0sEOPdTOr/356Dx
hEb/4mxXLH+HB0VAeeJAW/WSYNStqmsIcJGBx4lp5JjYjQ9krpHLixwpCp/8e0t5Qt7UyFBAefu+
P1PJdeyteMlRxZO5cKC1IelbMZxZF+qPVdQp9fWLbRUcS/fwrwxusjg6Jjl1Y6AAKrdWlFdv82Sa
Y7vApzm8N1xEFOaaGXS81sUuFRFJSbMKMzRfaWsO6JT3YGvqbaWDYTef6fbMsJ7czrJf8/G9iyWc
88PfOEIT8lkg9o1crr+Mmr26BZ+efAKzwH6ampgDC70RRvJ2Wh2yisrgHh7StWlXxtunDGAFRaGv
DZ83PKB50k0waue6d7RxXGdm9n6fInu4Qm119UjNYEVB0G0H3Y6cN1j/4wh5uX/+CsZd0plyntp5
f2cCPRNVBnmu652bbFalAD43j7LVB9sbDbaWPI5+Z7/9spnBOoIl2f8kXRT3Dr8qWM50Av7Z3qb2
zPXbMtTfUJiEto4e5LTzPEnRsQK8PD9Ewm49QB1WqsPssQdF9dSJY8Hy4Kphll3gQyKp58ZQhflm
EWHlymqXT8HQmGeIVaubFA/janBPHCZxUPU8cjLi8kuYRxI2vAn/A/Pr2luSeRPVjKRicn1TOrkZ
eKfS6lBuuBh9SXzK3kuafCrmY0Z62Dl2uyWe2BLJ9f0jx37fgZuGvkXEk/cgJ9rHbMO4LLrr7l8k
Ncl4LfBXk1sxL0F1pxo3/Oefb+v4y9uTuoloCCuxrGJsWO9X+SK4TFRvQDsqRi/mtaUHdPDGNZlS
DizpJPs4PCnYxcJ+jgGbHjJihdM5ueMi8mNFB5viaNYlu46Bpp2CFBB62H+FTj0/0IBUmgSisn8H
jrjFX35OlbpfWS1w7/DMuEyO8edsbQ1XOhNuWJBsEV0e5zvQtS1m8o7wGMo4cVuSt5MCUHZvhIP8
RbSV40YfElG3JrzvtAaFRsAylI1CDy9wUvAmykxxxljbefJLt1hWh3lrSk5d+YCorkdmtE5lZPtJ
WNkY+eP/+ghfldpPGSBvU+7B4lD6pOt9HwdKSQo7+qFPuMOPrIHbflKWtA1r1O2bJ8sINh3NmUQ/
AleOH17ZkZviE80wJGNaDwH+BX4s0LO8ls+cj/tZsnNyO34zU87/6IkrtR7Ec9BBOsk8ushoysWP
VO/VZ9i7/Fa1itmF3YlD/KyN5R1wQQcFbPRTU2XlefsDdgGzG32N95FD6pLsqSHWFxhZ6Zvy4ihQ
Yi9LDQXdUaBDKvVmN1bO0kJY6VKSjDPKcQQrPIsdGbzL1rNrSHlwj7z+FDmNeS/rXZMc349TY88h
XlPCbQcmPO2/SvPJX4jYSLyq7j+OdqnVSNdOj8fZ0I3u8M+HyEarGAPcUdtYULIZ4ZrjzGSMw3LB
3+KRW/jSyJwam1OA0oLAyyxBZ1NMIu7hzT/dGWxSMcyoofYe5Ax3IL/avhRg/oJ8yQw46+aiaB/p
NUSaK/Z33IDMHFrhMVy7P/1ksChwczLJX+tZyGrGrqdSfXH/tbaeP2AJI31ZBYmag3wQmsJq9x4n
oCMu8UHKIEMuCWl/8ObaS1+cANUU1O8LYv7vjWx0GiXUrYIyq6jBU8JwlGa6qZJi0JHSop806ee8
LDkszq/7ULUOszcq7D9pBJ1c/DNjiHwmlu8mFdDBoBVdycSJvlQNTjDUEDCs+n2Dk5+puWqLzki+
HYFnhwl+s+cI3jwLLx4kW7HyRf2/CWZtLhMXKxltzlV8wkqkuBQM8LLwT5cmHGhBUXNKC3wytYuF
AqnpF9kISzPMrWC3dCOqwJ4VQjrN/i5YxGKlMMEX8PM9ZIQ4qJ8vy+pOu6GXNqJCxOoehomtM+Ov
aeH9cWsO2ab9U2i35JaQDnPma+gz7o0UGkWRhGC8TLeoqjmfpUl+kRfp2lV3+BW7OundoerfRC9W
7yvZbFBeSilo8oYjnwPB/oIRRDCx87XYCQDu3WOp8Lg1nfqOXdpTTZ4d6RtC00owUiGKbWRyCaRg
FOLrLLJNf6WgFDFVHChNeqU0NXBbDUgdexuQ70GPQ9tvyhoQGTBjEZrM9NnukbCCMHy9O7sYmmML
tFqRVgLOs8TlWj+9lx7CnEeKbZK79HtDVpw3Yj80LJKDq3b+QALkKhpJNdExm0vtPj8bTUmCR9pJ
SDjXNl+6pusqVukDoKJzb49iiRLCFNYV2sY2PFztBDv4uazYxzJvLfsjSiC7dBiAG+FBQNwey2n5
/peRhx82gofegUqR5Glv4fvHCa9+wUFG4tvvEJ3sTCcgd8ftTaKVx7P8NVzmnNCZtbG2BMFsXObD
+z5PyUWjFoyDvxzq+elauElb/GXf099PmYG3yoM9iqkWq+1c3g/6wc0nqDV587+yGky2KAbT7Ux8
78FqK6SZQvdW6G3YSGo+S3b/gGlyfJCKy1PVgQ3hQoK7wakSVXqR6oVVbU/9JDtbjD3tNR6YouAP
uUejk7W3QfRE51Nxf8iOJgtyxXQBMHHwFz0j4Q9Q5cBIHhcnQbxfzStSOvs792UXlkJgLglTTJtC
IPAkrYOB4n+9oykvr2A23mj+0BqHAsCgfESVW+GCeFNJUNucYOz7eC+4XogmS3D37J4yrubPhK+f
U4k+Eam8Dt+Cy/78n3HlCXSgkDVnX+5fKReD7LV4Ru6O4dSajqzhIiTHHBptDm/ccKtMbR9pdF/f
JrZKOZayqZZFAVupRYehu080xk/zhX8QQ0kdLgyTUiXzcRCNgrlxhlGVt5ds7C1F6n0BIXu/+oFd
6FfCYjwXLmh456H21fcQ0yHp2Pd9FdR/zVBcZwoJFh63Sj94YOzzvhkaB6E1ZcysYLeeUVrcyvSK
IH0LuWExDH6VWo7ncALiP3hx/nTazTrUREHtJgVb5v86ZwQJUsZolxb0khSJOuxLlyQtylVB/D5r
PqC5CIG74tGF6Wbm3hYFChqM6nY4zUkMenLuq/uL5NBgDSScHA4YVlNr3NqvV4d8qrz6y9/kt/PS
TiW9l3HiklenL2AGLGyyrax7TvyfOlfrYlpgRNSOUQyMJ1MXCDDT/Pem+ekU+1wex4htsdH6tITG
ipm/IEw4DGcr1WIr4zC00ve/gZM4xIHmtT7WEYJoYaKmZ80M08JvfEJb3N7HJXlAHLF9AwDTGMbh
BXWVawbWdZW6mVfSCT25PeoDwcSu/bXhZTykkJ6GZz3XaR1mDhE0lIlb3Wx3Pftqplh08fVHt2rp
EfsTUPBiGl8AN2LjY6zglRYJCpA4JteM2Ud4MzHznjj8DlsPxjLY2LWD0y8TGkwsd3uY3184nuh7
xpqzVcOrOBL2eCcs/AwyCrmx9IAvquysDA7WjnA3JtDo+QsMe87KoOSWuitvEP7bNpcogWpilLPP
vAzerbbU+gTZbedBKLvx8mpIwjEuRTjdnVng1l+JFsTweXcWoBdqfiud087axhVXBy/w5lP4IPvy
r6/vL/xQP/oNtfthRP6PcTZvd0c8kk0K+rVVqBDwS5M6VB77bpKb1aIy9eorJHXlWrPG5gr562zo
ud9Vfp3r4YhaMHMldWDzthKKY4SPRZrCIaJ7EYQza4uPj0UIeYUxW0LwSuzj9oHwokebVANY8wix
+K2JuyngTG9K72ua2+lovJ5wKtF/GdaMO+pMgYcffHrpPfMXWdN2kOjtuU6nUvrYGvRLgEbxHqQJ
/0bIOSlFYUlzZQ94eU07xZ/DYKsvHozEDrdMu1oTKEKdsEJbuTD6cHy2nP8SaRfiqIlcImH9kbhN
yDNHPTQZWCO37b3LIpDZYvh7S40h2BxJUknA0Y344/ji2RpNA3s2Pl2aAI2iTYTjZbqvSP0PXPLs
2qtwK7eHRgA0kRg7nsLsSX1Rc3qH170vX7PlmgkpM02ibBaon0FNENxgsVHb8QphxOSwNoVC+JoK
xeh+wq3v8KXDO8lrUFVlPAweUpYmXaCL3R2urjBjxtW27SvU7Qjq8d3MSsMr4kl5skY1R7r4412J
nib0T9ViRN3jwlhjD0o17ApUPLIYJjuqVdpn8ECAGJ4Qf5HYDOTeK3doMZtklzVMiit5SGnfFmn2
sGMx2gZlo0m9tD8bTcYfvDaNiBlRGFTn4jjb95dGL0A0cg3sq9jK2NK8uUz1aQl1rBTz8fwVgpHU
nshx7WAk6dKAWWZrb4abU7ILGegdjrxeZM2s0wuMY73gfaC1ETCTseUzKz17srLmKv9JhrG6rLHl
g+BaE8mKiAxh6tT7GBvlDRPhIxY5wnWflutrKuBl9RldRq22XU4wysmFcneQ6vP+kBDwO5coiMKv
KSc4sbm2KXx78LGxdvhiVvTLTZL5zgN/fCv3nCrK237+FIdVSHd99g6Hk4K648JsBQPJGkD352GS
d+pg5IkWUjTy5+O7xZR7zu0+cFg69cLo0ZLPnzej28j0L1/0dDpt3z/qCdlZ00sswAeJKYnUjokJ
1b7tWxeE3w3x2Y7GX0rfb8GiC5re+cXY1j2tuZyPx9FA/GRN743jZBOkND7ye25++03wfkY1Bv9G
34lfFzceXch/fYsIr53In1S4FvdXj7dHV93q9LdzerasGPhmdZuzJRKNmyba0Cwux4exdUWjyc6U
dEWsOH12Wry0ISuEAbs9Xqc/pudNVN8isMaHzsikww2cBtRMZQWDGIg+f0oOzY7WjZJ+G9Px7fxX
d4OjFr5v+5K0t0wncVrWUsMJBGJhxncdUvpw4oyzYGRuE7C/phgS0l6gegXdP8PDzUC7qqcx7pa7
MEbkvrSkFCIIapqOzOMbQF3wvVxjBUUnIKbEoJy+OHSUiN6T1nfR/joRuB16w23vrqd2zSiaah4o
rdSS5gx8BGnfQQaLeXHIAst8KVVwbfH/3mNzr8aUS7QEPt5uPHuolyupONcSKvbbbnD+lFN0T39q
nZlURoTYJuiHwcp6BvMq0Hof8hoUl/FrjcpjKYpHjWcZWY53zj3HcKFhyRhmZzSUxrksdS3yVOQA
J2SUBKQgwcwDRTLtu5NhagfcRBJU/etiXxlRj6DAYX0xD5bkJTAm5TtxSc0tItFBYxhvLGifEeEJ
QQnzJIrvoBppfNP7WVz+vTSMf2jHWcYHfJJvV2MoioKeme1yxV3v/cJyFuvwFi+HZU15KEwI411a
8RyTSF2Z6sNXn3TyoH3MDoH2hmciSLpm6dykjgcvS0Juyvtww8po4p/1bu1rd2QWB0065vJXRcBN
fQF2+hLDpVE97UFxy2MNdYoH3CL9+I3gMceh9WOm3vnTbEYg/rCNimxSw/OvdmtB4Kvm7OxwZw+R
yW97/a4VjNVXMxYAJlhe9SzrssCUHQbUg49VTvOM6PrX7Ipv887zdHkKhfgGac70aSUtNtf9hvkX
nAKsp/6yvMNNpnCx8XSbgjUjvm2ZfrYwrg5nt0S9yipvFsOZod3JO4KXeRushjg06wpMh8xSNWEa
rtHpFBxUpSLtJhqPtAGAPnZgd2pMVVUi/lduj4hjK4CFIwcnumJLKPJ7thdTAk9upoGwUBWaKuxJ
AlexBW4dU4eI1wpi2QFrQr98RaTiqAYysTk8xt8mNUTyAo8L0O58STJ293med4crPHKEM44DO9CK
dorHTzOH8uU4JaJvDyOWmy9Kl8XANc275ZMfyKckbGSfTZCMKbPLSfA60xLE8lLeUkbQjQ7CJWT1
MYCpMs+XR65d++xZcqV1qQ9nc6sf6hhIJ0Mx1vFudr/xCwU/vH16SRRKbknccm8oFlfajFtLqelz
OSDaL2job/kDXjIq4w1VlVFIb0IeiuLIwuZCuI6y4NWcLY2JBkF8XnNrAyDHNTrf76o8lJllZ/aI
BsBbSvJJyo5RPu0r86oMRz88Hy0XXz/CuqSrb1bZJVcR4Pqw5YTq3Kag5LeMHdfxPJidJjwH0q/v
xRGd1yscNE0d0naXeafXXQozEN3RIsARB3ORLTa5RZwt7xjFtUYXaEW7Avn6sBJk5xIcf7/KWTJ6
O8flCS5Kr41cw6nkgQFChzPU4LACFvlbIR1Ru6koRG1/mLYbt4KELWDad4b6tVtsw++IFqvxYJpC
+U8tNFT+JHxyd/hPO1P+5shiHwFghoJ3LysQYW0qatsNl/HeLuEsqpzODHMqLeTEatpvF+HYimdF
SdVAZFMsyf+uoaQc3cnQKaKiXN2P2vuHUJGCHD9MnheZmzSScEkxRvtzf8ifhI5eESJhOQ69b82S
e3dm4q3OORxS34h+EVpU6EyMp0bcRmCBJVfjLTJJgy6QEzTOtbbS4f8QXsV8j/xzMaesLImM0ZMv
Vm/OwwE/CGbJiWAGWejZdJzMX0AbFlUEvKcJurrY/8GaUHLz+80QaqhITTuHWn6h3V7Df/YCLICO
f+OH4HvaiaIe9eQrkdGBcvYAsej3qo0sCBjd6DwAfUgkXRF63Hs0R1OTu3gX16wwNf9Kyc2aioVy
rsX7oAPwZ+HmS+5lgAroh7BC/MqBMmcoc2DdQ3dysU4yBBbutQKHtb6/a8NtXEG80tbolKbGXDnV
UOiEgeJO17mG4PsyBtqTC/niAMx2RDkgaOWxKmJncK5W0pNwexmZuJQCdfKJIG3NCVXUJqfUZFPr
7YOKd2rfmSRLq3eId5HYvHCeAFdz4Ugq5SOcJcOYu1INt99Q3I5nF3R40I1D2SgX5yOw8+urj1ZS
cdmPJKNqKdMtkn/6mVGQ3TuIphFSGMWn0Wx3VzoYTpBypvYeo7oQWWaAHVE8wBJkykjXvzAJCyc/
oXIRv8a92UaoNeN2pK8Bk437vJTWRJT0mw4t/BMW45FUpey5cQ4dhve1tpboWBvfCXP+vp1tNiaS
sBNAwBvnnpTwEXJGpOcFHWvcKCgjy8RQ2chxYlUBsFi/tEG3qPJRlTzZrufPpHeBFUj/oxqAXJik
Rib6VkNaCQfunHDUtxWbSTFMnpRI3cv7BqX5h93z78V9aC2by++yGTsmt2STw16rABBi+rqzEBE8
jcTtwWK6A/rXa1Y8dBJ+8j3qwna0UHBvmhSv2hqZmHL101sleibh9hkYWI/Q/BfNOWNwQ3z13xIV
yHYiCT5vPjbW76yqPBtTvOECHRlM+0juKHXhrgQh5duCdWjzhRP/ggmJrtlfz2aWsNWlt8ey0XSU
cp3MHJNQaF2Wz48dNbou7+115towi96UcdJNsH/Hweqap+XEU9DoEK03YDDaBlLnFhsoQw16Z6D6
Zn7n9xBTV2XPAD/SgPRoajG/yfPv9drtLBujd2EbJqrUQ0AwFZQss4bMRsChiUbl94dj+q/M55g2
WydzpgOyXHcLlYkczHbOxCgddZmlNHAnYwW909dpcXryMEHQ8+F2f45MVdpf2P5kpKielYb/0wlX
AmWVjICOz/RELRSrFhb/MhYIiXhOZK1KQw4uD4My2xezHhYW7/ZVqv9j+QKWd0YPK+R/icpZyCvz
8r6IbwvDZl2FqSgZN78MUZqddBf60lfd8Mwzz2qAupB6Sgc8YlaKpL9M8hxF9N7kXrgl3oirKuFL
GwSnAACz9pVQJ9YxVoPRUBYxt05OADN9VOQ61Z6S14XA5Zz5AIBz6e9FFwUENtM6+t7fDZtfRL47
3/GsRPCHwpC+xqIg9+/3jgSOuK+tCc6aH9CvaEjknkMHFPvJQ+4DrEWKksqLMlsxjNfs8xm+BLQx
TVFkYtePprIocwdvcSbbSDbVH/Vdk3rMCA1aF+9TbDbK3AYgaHFy7NVYLlWvcI67JTGf8Tx4dSpT
0+OUBq+Mdh8E1TvXZBltjorxmzhD18CByAQ2FKkBGReIxytV7VzilOxMJGnR6/WMpOa4LOQdMcC1
zcvnr1BvKiCrhsDEn0WuVIdVcj79WrkLI/9uapEhi7wmcG/uHPIkC4g+o027Sse0Rjwn7gkNtNx0
X5YEbK90SbROkJe73Xe0KPVao7MoJ03pqKHsOpIT0XMnPyAivSm3yELqH1Lj6IKz9j5eBWylf0Hh
0d6le4nSLJAu8DXmhQTfbFIPjCmn0ZaLojOyUiX3HOvquQKh05+Hoj10O9Cs9P92jsovB9tYuiId
vne/9eqntpW4pySiGtqaNv9D8m9kB5taZIGy7ww6wRSrI2+yPW2crHdzakBup961mWOwvW3Wt/GR
wd/YVBWvBqkwxggFF9wn1vNEeLmQBv58oZfrbWvtTqP/z7ONxa7+MlSjZ7I0eV4VIA13EW/g7JYN
s8oqLMgUWXEG0WZ6EgQOMevXhQuQIoRJWk1NUXj72txhmFFgwo4afHPeT4A7hh95IxdpkqKJ3nnu
si8f0IZ2H1mz9IWX5hqMKOHFu/3mtiac1ZjEbp164S8AufnilF1eEgBeWWYFvQiSYrOTErfDjjoz
1W+Z8QdYQN7LXVMjgZ9y6I6Sq2nGesnuEBLRqbI9WadHh3MHH35RyYdI9yzLKgleeB4FWnBBrnIS
SNsRFZRLJYiFhH1gFvb6HlOcRvl4Fi2N1KvNUbhU0kH23SpPsuEUMfhMo2hMdlRxU0dwfYOBVh10
pgqBk+35FE0NENXmCwUjas9llXJKrOKZUaum2pZaiUOGlacFa1tGuAasVMvoOxbpeA+TadiKxT78
I/0AB2gqN7LXhoKUEPvBhuY9icGX2vHE46aVAAO405vCOkwvYqUR4siHnmSFsVg8PmeDENDVpFs3
rgWOzBGC8sCEhNQdUQMEGZaVWRLlQrpdOogiVLTeGUP2FfiNvFBdyEpML/5SEA6G9DX/G94DWK3g
oxHvKH9rEKW3+8iO3z4JCcODKa8HvKUAfG3o2lyL161An4R3OvrZMIHy5+5MzATwXPQ6m73aVV0r
PO0T9a4ZMQ9GisWKmGY5wi0nmcyeplkvddVRVeHP66H6bmnB7r4h1YZQfA1IJsdFDwoPB5rt4JIL
c0trA5LGl77XQ38PgZPbNH0mxpT/wmtzi3riKPtxOa5vZt/8WemnjLIn0C/sIpXgxgFh8p4feUmH
D+aDc+KqWeWRPhTahuKwF1YP0r7untdh5fLYMq0y/SMQKn2fXZRvDInxqnO2RGyEDwVPvQwt9V77
reGVmvw3acDZ3IRz1rzitiXmpibIoFRsNaL9Ysfcs/rJv7hGDAf/BLINMtNwHjhdI+U12sICp0AL
hnXQXzYBr5it4KHjtCRsZqaCNO2WRGUQciHIkT0c5iXi2lUnBv87j4TbnJ5AdciouCqt+88W2mjC
iTmlRHK9KMEQXanBcx5VEmdQz3V1lHi6guE+LjrsCMZXTF9AYaJ7WH5WQpHT5JExk7RTD4PXIR6/
7gDp6Tu4WKFt70EABceExbb4B45n1aMTVLwqM6HDk8irv+kDGWdrjFi6ki0HhQSPpjntOqYWrAOE
3yWeKoZZeI62hdAy/21FuiTDgkIAyDrYb/MlMky75R4W8ZeYe/4Xm0N8HbQ6mKBHf23NgIewcLMz
Npui2DfHXbG7qmd9rPCq5Fsk9kflV5wRQO16Cc3Ch23D5sq/0ixRT9Am3ausDhIKqICfqyArT/1C
EwXhHeL/mlIBL3h6QxuMlS/Ei8scvi0S2TMDcB7brdFxGimMdXBCQUavuhOMDHQAmL6bVDfxCEix
Ktoynl2U9tK3BUjX+2khOnWN0u5j9FX/mIrbWO8RfFDgzgDPorM7y9/qbw37jnhQzG46zHEyrmyg
rLRAywhMeiE/EwJbjmF7KY7Ljfa9aSa1E5DVdJV6zlXfhAC/qPGeeu+yPdC8cAGgGZ+K9wdDm+AZ
6mME1UQc9/d/TUN7MOw9UBASZtMYeI3wFVpq6PJtuIMcId8gFpCD39qYPJw8gmznLUIzSxlBsU4j
OfQtEmT7tcTJ0wo6UJSWd7n3eugPTFAUoAz3ur1r1eWYDzRaq8cCnwUlc6Fox6l3JIKDsgqT2Cah
B8jUSdmvVMjyJ5J6dlFAvcRgdkSFO06CmH4qDJjk31gNsMi0ZtFyoJ2jf6MQ5eMeQbrKNR9mdirB
/oYfzx5bL4WXJoAytaVoacYqb0BjbVuPvXeTYRnFOTCNiWM1HO+w0iL65/YFzCSNXy3HZILsRiTF
sDEQD4ZL4QUFbq7HiJ5Cmm6g38hNvgDy0aHBMC3T0hasVMmeY0PHGvy4BrkBcCxeeW5tU7ijK4TC
IMyEg3nWQ3wu1/KI5SY2akOwOHUs22wkNlwbJGboRGGZGW7a2FLOkY4hyDeX3KC+RJupOLwNbxOr
KCTpX6VXtAbZ+M0YLsgtbSqlzKZKvNChjpMbATNOUNtCxMr1RwILx14ZgL8By37e2+TKqpuOBV6J
zulvBaTR6PMld7V2Q9nJ82VqIvZd6naV1IeUefTw5mlRkxhyGm3dPsSGmNQOSTm892vdweRFBIs7
kdJZZyUFJLIFA5iUPOg0We6RDT/RMY3pXSQdaiIkolhJ/CkJeeRmML63VPac7IMQZ+leGuQYt0Za
vERaHQ+ImWYcjd+4ug+WkAU41fgBzGGIGmNH2J1w3PRLRtObY69VdrrmdKN3uHZEviRyl5SaoO3o
wKt0AkcZ/Wf8/8/1esDFRQypkVdWrWOjojlABvI0v6o4tghMLGsHS7+oCY3CYZiV7LMzJPbkJhPs
5ASiTQH/i4ejEefJv7ZSnkEDd5jW95opS1EBTkfEnjaGkXsr12Ee+Zw+Lb2ZVr5TJ034M3hovKKV
uXjpQDrpxZGYa1hSi40+RL8wFvBDfGczEMGmZKrqNGX4cmZCbK86kD8GgHpLn7NvC3Pp4wppvTUc
CGRqaUVAOD81YHqoQLFumTq2PE8oa44Wn3iA6vChqIFU30//+lF/0jukqQbPfFOndTFJOIPUtRMk
InBzNH21WgnwgrL8UyCMlJTvp1hCNow5b4+3Pbiz3bxvJhlau0hSf5+5C/MFORR4C6aanaTjigCN
rwF36UOUKDV+k3Lzr1n1XEg/pW4o8S8P0QoF+D6ewjvmsbCrszZ6alwZkX7oNCWkH6pleRU+JQve
ft3WchUQaLqmt/hbPFrIvAgdUd/rambYdDKcmKxl11pro8OdYshXFFzpjjOLJt97Y6Qsi2e+jTGV
LamrsFKvz68ZMfmhfetO3WMG6PCY+08MxC3Mwu0wevdMfdtg3srUHXwIFwK4EIIQoT+jno0pwkbo
VKDNB65RspILWE0wcQSu162eRdAWbYuFBE8+oPkL0SweuF5OVgC82dVjphXbiEez4j8JHV3nfmLt
K0J+9qnUgMe90+GL1ddxmiEmjopZN/Lr3mdPYIAvlEp23Q6To1oU6zsFoI3Fj10IsrjathnpPBvb
wqiIR69X1uuuwq/C0NBrJRfcTaAOXjzDvJtztfOSgDoJPiDGsMYJfdOanXw0oSMRTwtiCwF7jGsn
ks+AY8aJ0qRjFTDvNYqU00xFH70TOopYTZ6wl17YOnKr+9vrCWEDBxq27/ImeA6R1Ykpf/aWDusE
srglmDWuWsE5oUKVcsXOBYGNeTtetbe7W5gYbRR0M5V8GP1oIzJUX5WQcd9BLozrF2I8Vi0ifvEl
H8hG46LZYccCDUyGsoE2G31KGB7E+VjEvktCJu2z/nIgXSx+FCxAz/xJsKFj3LhoNNMJYpa5TVxa
HlBcsIm3B/+aE97l/eanUwjHDGYr6FSgRfrbieWyO3gMHr6J15r1Q+g2FZODOowRElyKLOvs28Wd
OOAU8/lCvCh1u152CRTbi4BHbLTG99t1cUfHOXe06O++57P9KgsdL2AWYMITt4OlZyQ5Rovtctye
JotWEfZJo2kWPHiDELDcjrACSTkMA1CuqQUrC1Ta8+ZU4vRhc8tcHJF4dvqn4byPefaldEdb/kBF
Zlrj5fp2KY/RFVQjWUstyXjefYWbv4mL0o38WWne64ZHyB3YKpm0zQUJRNXNjv/EhWxtRq660Ud5
uuRZySKl/BI4+ADHY0J6Enl2t8FwrW9ZTq8Rl4eVFPkjmUwEhmMYuSJ8Nv9xbmsFwNQLus3n5dpM
auf76E6wo3Zjb+76tLAifi7vwi6YeUGqh9nthCFcihrvdwMvZsa0mj5FgZRvPHMGAl3W/UIzRoMT
y3rg4X30yogIkKQ6d7ib6hhmRkWXkFFCLWmQhN++zDx2A5+mea8VhrpwWSAoKSO+TBzLwkDRyxM5
CnvFDI/4d1npy1vRyLmhuWzv535WXTIzAdRdRzNdvkYg3AiZDXevrmabXzjKRT9H58S5g0el5v7D
gLlgVGsxwqAYR9SSueY2wTty3jqGUSWXwhAPZDBmAl5E0dH15C7GHYc8H2vht6AGAkestfIwBRi5
+wjQn0cjsEhCjKjMQ5L7Jyn/wWY9pI04BSpIZRoAcCmQmQ12H+MW67sTS3+XEsQt1Q2bfNcauy2u
axwkqM9OkTjIZ/hIY0s2nVKeC10NWD67MXP/bcsfW14Kn4fDaO+x+51cRvTpJsioL2R4B4tuOrr6
ilHsfd70rFqrA19SmpmVA8/UvwZlbUCu8DfLhKbBiVrnMdPwVnXSLighdimaWwOwiEgeqEQWy2uB
4I6M7ZQxbik14pxeZtUIKuNx0qkTitf2EUnD7vRn2DtJlairQtnxEjG48yjMp6Q8LL+q61Zd+EcX
kD4ENIUHaAl5O836lcHd9X9kQtBHjgdMMlXtktG8UaDb+6WIVPXoEKHVA8LXaBgfVEG9xrpHC97N
c1aAPF1PoU5JzIHQ9C7oCVV558J0by2F4GEBbnpnuzhPYMcyzu5DxWegjaBO0fwg0mq8F3fbqF6A
a2hTLnci8Q7p8OMaPXw1VPtfAjMOG6necz9O77KEjQoDt+ZHRy65yznqNRjJWAG5ClsQMSiJxOBt
pGfOk6yZUJXk9L0KnddlOwbHdQYkuExm8fQ3pYM6GvR1lQal3mIzw/1MI4ZY0ctU/+GPQSQoEW62
jNbcGDv0StubJShTiZ6qa9L/5Xj/yiucGe2PFMcBOWKs6IVR1QoQNIom1m/vAtGlbLHBGNtQZuAo
ZUi7JeK56g1rPB+wh07HS2ZuuJW0ZJR343qEePHEahjTUm573mGTzO/NJJxbTF/PB6ZXUsix+Qj1
uJTIXZbUqd1sKC2GqJiXxwBeIp+G2UdPL79M8tTAkNPXIETzruLWEkLjIJrwdDFz30LOt8MChmch
7kq/fIyRDzHdrkZiKku4Uln2Afd9cw+iHIOF6g/14rYIcctdbZfczryhm7VRPVci+uytig+O6Hzo
KN/THHu6Y4V30im3VBMyC7a1lTArWWSr3fcSFIW1tKLeXyFxIuIlMCsiXrEjRk7kzvpfjkvhIGse
UOLDlQbHAaqBTi1BbFoi1hnef/QN+hnzKG3Vr4pwpJZRySt9FigC0k4PZ/jI8Qt9bwtDE+wbfUTM
GASl9bv1Idv/DzcB7ZrkFG2ZvEvJ4ioist8X3627XHRdE4Kdm0a4/frmzAfD/xIHLex7hSMFpHKB
DXDABByw+aHnm7e3qB01QYCJ/h64n3EV1nFZ5rl5QjH+tiIRE8K6jsC2IInjwodRugcnC8SCCy6J
Db35UcbMQ/KE+Ur+J4Ix6xiCiyixd87lRgIVUZGAAKi0DXkKS5Qlq3Bp9vb39RZ8wB6r+Lyn1v18
lCFmUnNV5Uovo3KqczzOetjU87MW9OUWyuussu0hnIIk4HwyHRg7VvfgCOPyNRE/XrwS+AyfnQ1I
qIC/XviCpyqhOD2DlYT/8qBE40S/KGngydpeT5QIYx+EEFP4GtijDJVDfnTYvRY3UxLSRUEwKyBD
UgvrP9ZgcQgpsAxT6ZqrRNefFiyApBnmj6h1jqwXFUWy8Q1eJQTIa33J6CgA/CKhjKJ8szVOqCSd
mjLnrR4zeHYyCXyKZFQUZra/WN8lAalpMYlTPiFmt7bUk9MeWL+qf4uCadH7517zefCcW16ZI/xx
87GJyDk611CHH8zLTiICp06M5ypbvz85qYYh2metDSCP4+0xT8A/EwleS90u5c37sXJWHq66wElA
LkO9jhO42EJt0urdE2NV35VLKwqUh/kfh8y6Vn/HSsUCYDrcR4wI8xaQ6wzRqZYCWgsDejQwST9/
Ur1y2t0RQBPZWy3h9fD0M4VrfTjlrNoaHHQfaTlb4D4FHBLN2GschcP5MBmHZrgV7PJK71QkQEi/
9HEgpvpHf2DTRqVgoegj9+8CdJ2EA/CFnONPGbWeqyHeakbCSAoFFA27CKJzzt6EJ9Bdcw604jNK
chr4cvh+L+0eBZYWpYbu/OL/vHplE4FhlMuOyOaIfRDtX4vHJeB6m4hZ0R3LZL0O+EoY/Pkwsnzo
FCvoNGpzKqMfaCTkE2AdcgyXmTTW1GEtZxhd0G14mR0FUaYG0phXozFi+E1RPfpyGg1WUWX4BACv
pTr1TxdmI7g7mYPlzrzzc1Wb4FFF/gc3YDPy4lSrgic/GllCU30F+fQi8BTnYP3I+ltnaZz57bQ6
1vaZtL+/N6rc3EdIdylndc3scQBvxvctf9H3ced5yy4GEm3DuMWrvio9VQ3NU+9KTvXHEekq0+hm
FoJ1wnaleOZ7YFvOO73TMT2AOxTtyQrgs4XuuuDgxLXKT2gIjz62KTDXZrMIW0oKy2FWac+7kcq8
NFfWikwX8qrQMj1hT/ZjBiuZ37UZiCfPaJvJtvDGjoIIDJ8J25PJaYJh3M2zokURzDDukN2uvooa
f7lx+VFGvx+QivPOBVRCgMlUfPY55BqBc3Fly2l5sZa0+NGcyGZJmgO2enYOtdwrRxnWcVGHe521
wxZzbhpk+9l0AlFpbqBUZ2H33HwBP9A8Itxwk1UTq+M6hhdFM1sml7/zWwG2mrMdWUlO3t4voGyw
OnY59BUbvSojtC4XUD7Xx4WIYsmVjmncurA3JyWPGKlJWdFwOHbySJ0LcB/SKhGUYdWs5ZbmlePW
IAHkyeGZjtYywaiet9IQYRcraNILgwaf91/NkWivSAWSuc7QCl1+ZqaR5uoS7YWfZ0aUHq/6jikr
5YSb6IpXzew4qZi8f0q8RTnvDx1O5LTP0v32CEXGGYSUsV1vqpoWRW7O7pPyF5eM1g6A04O1JZhw
VP/WiUAH8n6DD1x/JogR681386rm5+igYzj6farurBjWSW2ALlE0V47iiVH6i/VOyNtDrSEa27yt
I1vcfaAgW/BEEkLFPRV7wUhtznAII/K5ucaK05E13i7fTo/WEJEwdtimAZSzGSck2d5FGh+otU/8
cYeEKiO41WzaBENEE+MN4ASCWDf0zWAejr1qB5ED7PJTHF/RunimbB4dN89uaO29JIcaVHzM1d+I
DXVNudIaY2rK3mr+oIwQFCh4IMdLsggkHUiCds5NFKSRN3i85wX4Ps11hwmulsWZikfGiuAKnpGa
yiPV2mquXw2PqN6CiPsbvvkbPnBJn5yc3bVGaqe/q6+o8WShdTeSScCpoxF2T6ixZbycfKYX1LXj
v4ztDFDyiyjI9S6Kd6JjHFjAcCgqOFATF4fumCtwL/jkkCTUlKiqml8s0776wcq5TssSXgYxcON1
zukx4GmCA6I4GMnE2jkZ8Late9uIrsyZmFDxAcb3IPXcxkj7vlW3XEzfIZVX9wzR9A9AVrPYYGjH
6Q2ffbqqtJ5BRQM0Cfp/nJx0AFYYplMsa7in9N85Std02ytELDZqr6upmsGzRar0bbSro4sy2MU3
rmRE/F1dr0kkpm6/pc/tftymIdkJ2IpTUUYZ6pu6WPh/eD7y3505IXUNBjAUR9Ni/xRUHLqzTq2S
F+F32etzVaWIQjxzzxfG30gIs9D17NiJrN3Vw57QepX3htaGk6t7hp+jVcWts64OIDFM8oyS5Z/z
rCJnlJI8Eb7xvU3b66031UHF6RaJ4WlbLHGFid+rPTVhzItid/KtZ+BzhRSppsjDJ4/79hAgtsyf
Z9FZZgRGN6OK8+poVC6yszCrzbhOdngCXzmia+XUxLWA+9nXT+I8pU3yJKxmTJ76jP1O73jLbeVm
SN9dxTBUsdPYetbFUcjZPTxrk29qdRAT4zBYRJqIwvkAEB7TwFbT27AXUlhkjrxoM5oUjZje4XBs
adphCs+RMMDDDB1pNx8ptTAW3gp3q2UCsK1pGOXbai3bNT4w7kEtWgzaVBAiDbojdgqGTIZMskk7
4++sGWKxWky+0QFFYcWeHn09VE8MdKNTdMpDgOobu1qylOE49x5u19qm+AWYMw3YsU8CPM1g+Seo
Q5vm35XNW13pMPWfgJuSMoG8WUXOJ4JMqqxtINatzus8PQkcHuVtV++jmqDDa/szznUNL/tQdgJL
PISBPqYFpWBB3ONFRbrnfDQtzVOP3tHRZHE336rzaAm/9Tyq5MQ0NBlyf/LoKlDWG03wajGiDdsw
sp1+oFWYsvnTnJ1Hn3gfMnbTuLAXG78EFBxngPWrQVkDtkCRzIm7aZdMVra5AugCin/mxbHKj/RD
6Zqho/DWEThE/Wp9QAI18mEghJx+4ODT7YGO8rurQukwKRJGuNQYPkuv3BF93QTt5c+FgLmmIOtc
2ME34DSaeo8d2pA/o26rP0oDTeBn6iU8zGRsifcghr248zx/5KbqE4dznuNsoU5hyd7JEqS709kA
+iUKAJTifPj4qLSZ6HhhcZeutNxC8TSOtbBfwnQ2nxBiyuXMhD+zz+jK5hc8zSR10Uax5l9dAV1A
9saHlZjKt/+vXfqz1Ce6FCgR4fanjJMhGTl27ZxPDk++zZ+QXACXuPCXXbrVtJ2JWBhvZZ6rzz/0
UswBEP6ai4nmaXHAplZ6YmgfUuPXUede0uCywxG72DqefGjyea6MRf45calBpbgjypXkRt5LMitO
8n8hyz6IeOmVSmMqQJj0xMb18F9gzhDvIdhx2GXC9RkTKI0vw+SIOr7GEpn1c84Iz9cC0H+KurC/
cya+0BNSjgv+poUKKxo9FLxWUYJb/PGRVyjznsJ1rDJH9ECmhyD4UcylQsB6DqR6Q6Db0GvuQHdL
2Gba9xfuo7NqemVwz554h7hxFm+8fZ/U7ex2JjEuzkkekFEpQD4BHPkaY7yrb6ZVFb+eMYj0f11P
UFmx81lQ4RDMupYmVvJHnLXqZC2dFHq4KZcldzt28ypHhBP/kqxjZDB6HC4NVdm2xSAQUaYZoggA
c8jN4hkfpd6EJC+j1TnnaZ/e7AoTxzzxqKie9KgLY32vRSkGRbJ67prNfOkHWd4gBksyhFnNsBgE
Q8BuivsGzHDrsTPA3fdPb5rIe+JoSFluhY2wDwqWTKt/eXtqCmnvVX26S2SWZ+rxFZjCn6JLrt7s
IlZncPrQISuvHsGeN6i9QUdSKOuampUAQTlh7Whtpr2XcIS6SPr5ERyztl/yorl5DLPqgcvvewVq
2+FyPp7uK6/onQ3PfPPq6mXMaz/14o5fQtAM3J8AitpcIpkem9B8tfbThrX4wh+zGByK4yOMzHJj
h9EVuZ/b/xRUV3a6cQ7siK8lv8RrsIhAi+nklgrqafbEgczBFoRa7YIoWMM9im/K/0MVqUXbbxnA
0VIfffnfpi5XbSM36K2Ijbb1AiDte+5ELhgFRnJ1lveZc5nMPzj0R9DvLgBLxj8YbK2P9Kku+5+R
iX3f5fVXfERRVRLe49J3fOqsJTfoxzs4uPnjh/CInqoieYrDyCRETyAGwL/paP+AN780p+R+t+Mi
zTiCVQU2PYNGRW5FntsscZbZPACSqOIPVOpAHtyOpX3nxgOtVzqocctje9HjANygH23DXL85PGBr
VY5LlCVMmWI+vd391e2No6VcTQlriRL2RNBR2wx6i0SiitrVrCFHRKDQgTniYYNIg8cxNQZCiAo9
U2fIUtjmVokq3zUf+e/Mx3mcJ8E/hf4e/kZ2afiKMKV0eT0fxvyEOux3whkvrlgSoz9qXwaxOIG4
6bjxnZWqLLb/SgOoom39VEXT4gZ1DxRdwgrbo7ON0ZkiHTFQWQhzVvk67XuSkWoHbr2JOLi+cz2J
dzAbidQ/cd8tl60YzuCxykhs3R90DThEMPAWfYZMHtskxcaoWFv2+BjVFBQO6BOZbNvmJ5MhmPdQ
jtQqG2oYJZXH50uNz1bWPauf2F4HkH0apodTte3Y1m5jYm5dPzfrXjycfKzrp/8UshayiuQwYl1/
0rFUIzZ2gz7+UHIMNICAscU57RmleGiRbZxyx9tecO/PkBVJJXlSLX5Z51nT/PB1DK8JgPRrhv/e
tvPQJfxIuWvrYcjEqwGZ3qMR/mgGZQJggTwdiUjE6l1OcmPsJfUOB7qGNwuyJpUqsV2mD6ziegLY
E5E8gzz3xwPGzUkZctRiX7reYKx4Zw6RAJY3wJNvvhqzPmrsFtoAnnvBX7vB+4V/fiv3EK4+xQT+
8bB6DCr3dPT/RoET/6swKD98kn6cNogaWzK5BVtXgp9/zdqM1S5dYfs1Unqc7DDWu1l11DzW+qVn
EiqQUsly6DGfcpfJzAkZUbkpwE8FB36uFF1k6cyLH3jUIZyqoL1JjEgPAbrFhLf7d0NuRnyr7yqD
54Nm2pKpBbRe2avlAYjb3qaC7t3IUEyijUBzejEVyOFJCTFj6nqrgzTzQwAbsgWIjW2dmGL9VXzq
YAuHuGHXXpg5FvTjC8r8ruwVQcN5BbJ7Gfy1HhT4nlNTssSY9e90bEEHpjBNBJNMg5hzte2sh2T0
17Fw6SJnQWEiZddAgSJHpdtVzoDIKRqNdtk39bkhFJnrhqgzUGcYb3oM4ew1jcpCXGUL6Xl5hQ+u
oX/2xSUFGBlQ+buAO6uA0uRa4jzlczvkoU19sAxfab3Y2g1GH8ECtDyB/9ESTll7RX8MTK0iwF3v
Z/s/PKiOGfWePi19shzUE9lmIK4dHqGbNXZeI+ycdxcs+pV+ar3gdjR3dbiiRMS7zA7rbqbGLYBg
Pp23WLnH9AAdghyI8xOoAGLNDeLPfOU5PVMbWUKDuy6DkQWiXzmoIHoWNqq+8gy5XoLmlD4oiftB
ifJdenKJ219l9zgmCg+vHRV7bs9Gw7nuOl7yC2DDC6Cut9vBOTih8KZlHdzvdKpI2ho6Vq0TiY+x
QMry7WiiUURU4d9YGtwCs/SuwEAh0L7s3RvfnW0o/2nFkqBDqYV5jSvzCtu1JTZhLb3EDygtCaWD
hVrhzOdEdls9Ov75+/m3SXW14FkOFqXpxZHFKfj8jdRVabAK588y9NhKu+AvLEu3gwr2AUsEvHfv
Cmh3kHdx7K9+O0QatCOCY3ZTimKehlPoASOVA1Iu1D5apMF6QV7q/ROykZ93kKbPvbIxJ8jYlsik
TygcfC7PD4sIF+QVqhK6eEg7ABVDEMMlfNZ24FsszmS62NLp+LMcz5wm4ySWplfc5n0VVKiU+45e
MqMwK0x+sOCPJUmA6THAFhsV6nM5Vay53nKnN2UpcSAhdd/XPmjEpIkdgQji7GR2vcMuYLhA3vE6
j3BCwmJfbn2RlbZmYa/rckKTwB2bo/GXwF1g+yiJltzWa5PNenP9RFkEKzmRCbkNNdSjbUOtsnqF
f+GtSb+rb1vFU9m8rDsXJeJcz1l0nWoGWU0F2jXI88jrjYCMrfTmiF/hCPGhXIb5iNU9khkm1PWK
kXkLgzxvwlfsGHA4lK4p8qtJs+DMQ3z26QFHFycFRcIKycP+cS4F1A7rDxsfx6FvF46EQjGRLUy7
Pfem4s8k9tP/yxhIkWsIE1ieGpio8y6Nun82TLEPia1fGqaYghM/IKGKhuS/vEk8yYZh72RcJUhf
XeS9/39FoLgaKaAGJD+ocL+RWt5vGl5foGU1pjKs9BzMss6RYa/azutcWUtEDaZpupDfuL16n6W3
yPBcZ5VFufzl52joBcv9luV6OKbCifiMyh50QsIIscfOJaH2WsfvapkfvJMt5BPb9OgjsSkRHzNC
nSinRUvV3HxYMwlVn8GuoJVelX89ozSw6t9+kL4M/EtxwV+BzW4KqJdSbhKxvjbyFRXQzh0EGFCY
WmFTmNi20jFAruzRAWTRgZGZwg17dxaJnw829/q3aE84HvjNP8G8ZlsRFZcIwCAf1WDyaXO4Mmq0
8w08jTV+7shkmAtXyrMOTET5xxn5cyimtU2BX75JSB+IfJmCtLmGJnOTZB1TPuQRD8AqtTvW7uDu
SXk/179SqLzrBfhbjjnd5EMdmd1RnoRlmiHjImmwTFvkwZm5p3m458NQ+XODkiL3BSRzjptR65Do
wOKOKiuz3zii/ROztHNMRK5B4PsW77WuxrTzDI6HRZIsgJ0j52c1skOpX9nTm1yPnFIBVUWoaScv
3LzffK+dM6jeEWpobmy3mAMKMZ8xAPKuZMU+JCionDnTjp7gAScJFLPcs0Wxz6Y0MTlXjP7MeOit
em1m44OHVsJ4BclMFOI732chcKgihanf4bjzwwc9vmubRoa5sG6ii5gTCvp3+rzR/WPlfk20hm92
txfqqUuFPABbwrhMN2p7P1y9Qnv6EREulEG1KgETxECx11LIO/S1g2m/3jXLJsAo6yHSsVlJwM4j
dJWWpFcAdDHNl/ukXhzoN+je7nWuzbj1IIpH3aVCPfqp8JjzaStkfiVxBMbH8sHVtYzNDMM3KHhc
SpcJnZNYx+reKly9NpITjYssElzkXJ/HZxe+5uqOZMjUqTDdEoFbkiJ/85/gBmXut/kS5QlsR0d0
k+dnrk7cQn5ePYw212IKwFuOzlTCv8v1Mrero2ylskl5VCEhCFzISyAhomj5FdQI6WZwsjQrI0nN
MLBHOmf7gHCUdwNOI3ZH3S2zqR/dpR481nMCVJcW1dVCqe0Mjf+LkDw6rOGwAMd6r5+EkrxBvdDp
kvB1ESFHeSbyj4h3iRT4plNp7/56nOysS1BsB2UQdEPRIvnQ9iVctJRcxp4rB8DlChCylQWyOims
8CrckSCeM0dbPtxb3YRL0m+ER7A5DbJB8VxXlAgPcVdOJOakHcTLI0vjvJte0AkuPNlhEaVhz+8s
B8er/6lUylv0HGpPB0d5QW5T95YMCIWebhB8ovbx2i7ek68UMhAitlDYsDNW/P0bq+2/RYm4zSxZ
QmgTH+XE51K4ZRv8iMedYnGX6x5ii+QOdLIwCmVy5EM2hb/+wgKw8blhkUM4VtTg/rX5LY6wkViy
CfFmXcp1YOeM3/KYasbL+qJyHvuLh1gn1DZUEkJLuztoIJmumQbTjZRqmZe0ZL/YAaCVrTWWivYS
wItBGzLISAstpQFDR5UUlgucqnij5CC5kk1l26K0QOVEwFZbPC5Proykr0A4i6IoEsX4YQBfUtAF
iG0ncCblGzA62VVcWpocymtWrAxqI3C+KbQ6jsm7v1VOH6oQD3xuT1a/qqUOQce9c11GVTe7ryJT
jU2Rb14GMaizDEL7pNUHaTRq7JHBWXBJ/OgQSGMyamvZX4qsmDhmpH3d5+T89XMWqGnWikpf3yOT
iPFfWkkdym2ELAMXrrcLpwHinoEEjSOqhJydUa4ZusaxWa2TP6GYc7Ty5fwIs7qVEZBnH/CUECqB
XHWN7XE7K59wJiV8KX+jGQxgFqm8CzbmSpApAKDg5qXR6Wped2mhBK95+g9Wka582zJiT/sOzsl4
6lS3Gz/KMvVk4FCzBPIwT/cWnayi1Xv4txRvi286M1g1IDJPjVNvErudP9Cn7z6jz/KTQnK9NcbE
0JsXGz5u01mL/a0J1dmZRMDF8in0ZgINF3EI28flQfiP4V7+ySFemsKMVhF4CMV8kL9WtGaXdkGh
duMFXsP1Shh0avz+I+gu8jIu2pcUEfeHqtIMZpdVuLq7O17n75/08PSJtZgR4qTfRn3QUHEKomId
D6erAMEl6zHhcZnVAKaHq8Gla7YqkX9PIC9G0ZxQGZSzpYbAzd9DJNNN+XQFlDtWnBq3Pt1lbAwq
5YL3sLj6DFbK2wPPUwjxOwdI6BJNEZy5VKFYyis+gG0ZsRnRReXcCUtN0JkJJXYU8NsJ5n41NMJD
Gky8B0eONrBib0eTsvmC6LZy37KwyQiFIz5PfG3NsJ+6nqhwYcQHiOLgsx8v4BxQPvu3eonN3sNz
1WCkW6hkYiRwo/uBlMBqm8z3OOwncwSoRdKxfD/IXD6ZBhgY79ZFRHuBnqhVWxRk0wTLi/zARZWp
D2H8BO4PrapVSl4lwUdqyDzmQWgWYdXsRX4o9KgsYGF8Te/iAtQ6nKChFLO7xAMpeRwc+//KKOSo
5mZ4chHp1PEYC40tNlN/InEe71SV4ZPl/HP/x9MhOZKQf8yZmnptZ9GaWb/IIZPzvBL9U0refQLO
+zhyhiyf3ZhkwgCXKlJfBIpUZJ/oFMBKIIq5IJ1C+Bos4FvD2/GX5EXxcj4Vbq4wv4EJd7os+zGG
QanDrkRZDMveabq8sWGDWJ0CMPcxARh24whSWYhLs7nT69vzemRWtg8QvSfjJ7B0aYHTDHThyS1D
zwYsOrCgknz7T3ffSWvfVjLUfNDuIuxc+mQIX5F/Lacksj0wG3JKggDsrOytnfFT2m0Ujz0LRX2m
cBuwlM/bFQ8ahmeYusjSCFVb4WWUa+qSUg6NFqHjQvr+xYdELZBa44sJYqOYyrNVGKsKLWqb6/mG
B8D2UulSLxx3Ha6Tnbvbs+x/Q0myD5nD/VsWtCZdWjVKzKnwxzjlLXyYnSNm1d4JqMD9Yo8Ph065
e5Oxbrhc/eII+rzuSU8hBDc5q8yiIjt927np3i5D5VjvK9ZexEG6KVS3+M8jYcG3bE9mwYq+bsZC
IW17HOqyE/nK+ndNzH+F91wBL1B/uDhvyj5T8zaAM3DEEFXFN0Jen69yBj5zUoruO6r9LsWsOoYm
Hm8Pz14oRWsbtll9zVoNSy+Zbb2fYsVcDWY70Y/7Sq0iVEl8LpyBMKMwjLN7uHvKs+qC6ZkaPnqt
F302b4Em6vfjGkwM9If+4TWBN8e8OncqTDxHHzLHlxF9JZorK10b3aXvnBHxZo+BtDdkn8C3fJSZ
1A1qJpjDYBIL30bskZCuSvKow0qLclkScPkn8IgsMCF+m1mQdQNTrupf4/l374VCoMQXVAnQ2V3H
3+cZbNi6wuIZO3ztkOYsTaaTIv+PZIIMRW2ky5iaT56f2EiVtRtuB4GoZNMDOZPoPqQ8ZH9zDOyz
CbTmY5Ga+yohYZYLU4gB6F+ShJ9UUsBdaFpaWmQN4DNuPw7RYyWFEClpRyIR6BQp2OzmZVeJ6Gqg
4g+VtxzA4zJeh5hoVqlHnJQ9GndaY/uZfqEZ+nNwJnYbtLyJ7QgJpbqQGJGZv5HyUGSCIReMCRqq
iShRFhie3qL6t0R7Ami29B9kzCa3H9vdArX7rxzuZEDT1lsNRrMF2BaIWnetwF6hWbHNkUrmoH+w
Ryraw1UDQIhELt2DGgnWRES34kGdnI8sEkSAWRKZ0uoGzcf/BpftCX7ezhz4+30lgeNEBZVhiqTq
IO8LzbYV41cBTp7HSWQBujgehYWMe6nZjcJi0JXUCWZ6BABI/cDgsN1+ofml5PSJ0gu00A/x5f4d
VjgsuPyFe2mwDGlEvSMRBarrQQNIfBASCU1hUIzmO1QUDcGKPPbaNs7r9lO9iBsnnS2q24xCH6HW
xerkorlHTKSdWuAxsCTjW+AOY+31u0Wcon0KOuzU6liUlrrBxNH/TjvyazkZJt10fBQblnJ0x4L6
ANEQXZLQiUfuHSJHzLGa3IxfdxKnAUhY0owvkwm1Wr8lUvnfgug/gUQs8zRNFGiJ3ks2p84dqclB
N1tLiuTYBBcv7JpyRXvPwNK9CqYhlW1lIpbiVKR1sP0waCk4/15TJokf7fb9IDbB2OeXz5EH8bh6
hI7NdOfEml7YYhVW6azYWi2AkhRNdFpqEvxTsRQyAv6lODatlPOKNsdCbukMEKbvbFAiXJR4I5Vq
ulxYh1FlhxLSZbi4cU1n51ibcBs/1YqeS4qfExfqKhw6pn+Ef+dsO1zeZziNtda1EQK+QGqya6l4
QjlM7bGixYMP/oD5seID2bt7NT3e1HWfIKkA1B76cZehYmym3mg+5pHAKbA92+YPiELa1oG+guvR
GVhosNnoD0Kk6N1gnudR7W2Q+6Zl5IfhNOwQEZItYxtuUXHW+ha2ilMrxb/dDvkGRDaHRgT0DYNO
HRpi6Q/W0gyrKIcq1KYqJ4nGyq3s/GYnK+jrz+f67yeeQqVojF+9/U9Lwt2lGSwV8PL0Kikg3FRg
trNOPlbhgViHsrCeHIz0b2B33xwp6fm0x+C3YXTUn1uLbgZ3o7UDWUA4+QPUJlUXVvICWN9lp1W2
bYBJu4J2ZeLxy49LiZ3Y1CTCWIIF9HgMHkQNsULW1YLy6lJHk5Tk01YqSs/7vbwe32NsIPUWCZmE
nae2AEl/DYx5JW0Pek+6/TfBfMnJbHV9pEuz6p2ZDVM1T6aQpfqdip4mgXzbEK0kQ90pC7Et5yze
WuateuN/BMdDr4fye7L3zsdsUm9lTo4z0yo3XhM43wHgwcGubREJMyi4B9yLpeQC+iTkIVKKWUiq
Wn5Ofau/JgBmPqkOVrCAnlvQ+cT/nvkVLwSy4f+hBVmLtQ3eo5+6A/IiDjRlWxCgEgXxmOur/D1q
ymnuBLOEkqcP/JCc2FHbovv9vFO0ZRmh5NRiZdpnxWGHlu/IOv6aApWyiXN76cX6nVSoVLRJ4CY1
oa8TGaTmkZVtUrexwunLdFZPOq2Hgy4ef04pE21GnRQQYRUXVGWng86x9t123jzzgA07XFaLQ3Aw
keNjpXMPjsJK+PE92GNXWxNzT5QtpM9Z/mOFpk9IllghV5V2RsPWbFthwGftJWdIGK4INnPE+YDX
o94M4McGyiUeGzVPWTzf5s6H0W5J/2KZqwLUmPPclwxHNDu4oE1uE6jgp7jZXjPEQSieO6RKo93y
PXXJLpZb9fy7amXcRuDpghKaSJFHLr6kYQzfDKgAZshm2AKVKQB6mg33KdbjplSIm7+2TTGxsVFj
XQI5FM0ARf9IA+e1tBcpVFTeXx39xYcNoZm7/qWJfmkfFuc5k3BVzEEQ1S0QIOkmIgI5YbIyo0yf
zzaNwPioSkaOrJpe0t6rgHO+3OlUUSQWaLn+IET0UX7nJXtvjdTy3tR+FrPSkeDzVncJIg2mz5UB
zhSTugcPJ8xGVwTQdtscM168OGOMW8n4Lsx25riUQNQr1fsIS8WRKcQ0V5zWJworU7CIE9SKaYK2
jUdcRyx264tEwESAC3NXghxO+C2+uGEGBNPJVakld7eL22PFqa+q+1hScz9np+ZE82VXXAzYl2i1
+zbB5ZHM8BfR2AODQIO2CayH2QjNp59AIVGxj3T1ri9W3RLuS9Cgvf0MFw0byrM7HDxNl5XbnLGH
TwL/GGfgseDWvN5/Q+HEeC1w1IDibig8CsyBZxJ8yOwwk9CRei/nIZTwUr+xcIBQWNNwlYcKTY+A
SWsZc/LIrLzrsYK3ONZXHb4yIxln1TQhrvWj3BcybvsekIFAiyT48ZI21UBPqsgiAaF87YvdLif1
+cwwlWG9Bwg8p2RwVqU/m+vOR+VFsMJC/TcC4ZaAF0bWGjtjguY1QYa33nV1NA7Wd4LQ2RrvNMTg
Py6QL4L23BR/blnxmlWosQaXas3FlDsJsa1vVv4hXQj492OhU84+vMkaf7o0wtjvr2BU+7oHB4zR
RYTlFV//OUib8r5dqp+IeB4roiEEfPa2QTYS2oLSE5Ixsp5r68DkCHzApXxHy8ejO7Wjtpmtplp/
xTkhybgH0/WL8GpJKObdZt5pbMi+qq24P+Q1rN/IlQyBNHl6u/57CoGLBkoG/Ii1pdwLKeXrv+3L
P9+AKWBv5+BL5yh4j74ZhtW77CfNDCL16iLhLztvoTL1qGmKGVy9Rc7pIE+EVDEaf/fhGKVjrfig
6kFz4XBy3+6y8I0vROKMSbOHdlGBM0Rpfl+3DkWwUnuCbb6udQ7JnzbQZMdwv06V6WBFpW0gdsWd
A5i0nwA4Av5SLPyAEOLi7/R3z6sAAgHd9ZEUb6C65jdWX5PaVm3N8llXevbTVAxpahc7CVa8gufN
dF+vdkjkHkz+M02wUTnuZ9/i1yOju5mwQIzfL96iPo5SjHyF6g6YMEmpFRThnt+hkoIed28hSjgP
F7Z5u6WD4TTlQQloTX8fky4USuWkC3d2dxA0bXw81IYiXFo+egv9xIDM3G1gbcF1hI0ruEW627Ex
rEVdoSzIPJAJQUtmtXjkJiLMu+beQhGasrPkAGfByGlq3G+OrU7yEoQLDpnUFfLJ83Bas5GvwuOu
n212rumkJ1cyN0pMN7ufx3JETGaFlMeyMA17WdNpiRAnLY7Ik5SEOaMbutkuCNpLpLno1nKFWtC/
5XyBzztYXJ7mBQTrRpvAp//Wrvjoh9f0p+FMx7KpfhJrH7TpBPizFuiPH7w/aMMfa5Kh8RryRa0n
2vUrbuadcd/tX0j9LpxUb9VxrDO7GEpHh1M+dDW8DdBeR3ARLvoHJcGGA3dX05EZaJQtHG5pebpd
WJHC1UTTfjnRNR4TYYkeAbmGRWHw5dXUSbJWr4wzCRMOabtmNYcpI0QYg9NlTAiYHdi+EoOzlN49
UDuMPxur9mOBUdwp/McEnIkABQ/E298/DhGbaIwj5z4HcmQ8FMULyTOJLWP0kKMkdhOV3y3BvbhS
L5G4dNea4NdM6/NMmLqx8l0gfkoYPDtgCYFsMcp9AtsYcoQvH+cxQC0jndYRrqQ8jY/owbeaN/Lv
c84k+4rL6M4vhGSbhHAf2Fjb4NLWNr/vJnMaFpsQbiLePQFNKZ24USuKKY+IgFJ4EEFCd3njjxoS
1ItQJLkRql+m/eYxzuF6MJ3nlWc0uE+FELazTZfvauXduMk4FSfkIPkuzzNaQfOeKTn9GytNKQYo
VXMGXntDv7GV9Giq6wRXgHCQHGJnR/vXV35i1l2MfQte42gDCrgT0yYAw4LKZ7F4f8YKEG+28pya
KrnDHnPgdGHGGSpwnHvWAILrqNS3NB2gkwcmKu5iMDFXGMVOXAYTmOn3+qEUJwzDTU3jGGOb04YB
t66S4NP/oETaTEW/gyAN+kmbxSqeX/+D7wyNo5S6DPHlXlxM1UzMWXux4tgLJR/vjJpWro+kuFw4
SrGJc08rgjU5MhvcDftrajzsvYkm+ch6dj98HS1a44LkZ5nkB5akBJcEDxDd/5ka4RHxyQF+ThH3
dG4z0WQtQaXEFLkyW9pLua+gN2musZ4ulCLAlM00BUFcmo0Yiv/1oWKJax0+iNeBRRaXp0z0BnkA
MHQR5pDEHTvuOeQLL+yM8xoPhVDffNMUs3zxrBzXqwtRsjhx5Ni7du3tSDMTsgD64nrU87wEDf+N
04e0R+YeF6p+9sVqVF62k4nsx7a0G72ztpXBe4MmMHUyJoUtxXlUlDOFKa6ctVrQqZURJ/b7haby
X6NGvSZq+LUo6eCi9LI9pT1zmub9P7H72MvO6VtBUX9jS/Q+NFB3/XP/cYBByJ7qOX2vhFNGf0jb
Li4uZPYCW3thth5BKhR+wrkNcrQLv4uQeqth4QRFbdUtPCTT7Vpyqm6za4BvNTQZDBQvF+8jATkU
bRZjHcSJjtpwyF+WWE1WnKjSlP76ATbHoihp4jgsWOOKfNh3dOy+j8+ycl+fgl+Yhq2sA7/ov3JG
kO6V+HSq7icEyTSAiaDT0wogVjU90kZIrz4tD/jAMSiTAArjkVdOsgj+8z5SJHKXbo7i4AjpSOjZ
HfN/3eDZOa+kOlP5wrS2+BadvSaNxQi8/T70B2tYXFzxTmqKgIfghM7a4LZ5VoVQralqeCqQ1ITn
vXPrBvdnugiLrxRTEjS281QRV8DAPlRgfjEzcd2hWR8RYkcm1xE+pLGejX2/FLCdzl52pQMkP2n9
gjS5pWjq4AhvkyGAFGTVACysLVscgo9WnCk+1Nxnf+WMK/miad2McDYAfRW8k70Q6cNRV9cGE3/J
bscNPeiVDFWf5Hgqc1ptPp8Fzyc7XN7uP6xcm0neP8LlnYbpeqf6y8gl+pEV65a6FxtG1WeMfabW
aNTWYNm0daOchBzJt2T1jL/zuEXTXsMwuh8L08aKDv9HsWHmW+v9S3JNIhMjXX33eHtBWA7TQCBG
Fppmsrh/VwhmAKG0axzDc3crJm4kH//qjWC1yBvWZLr2v7I7FQMrXA+kMMkbui9UCo032Dv0HK4i
v1Dyjogvd+yXHxyfE9ezhQKG8tLNsHYWGKUPb/8CcK2WvRqajjAlqUWRX8z3Hzha89VblClRK4Iw
yYtNGn96Z75Z1dFfo7/qywywh++hHZcziIYE8qttIaFonEWx1G7WCm4eNEssyG3aEZkJUKicV+0b
DZPedr5QwfWmuFbGl3LCmaYzFV7yCtDLCqO9Zkup7ddWINpZpPHIu2L7tsbfeMyKlbiuicMQeDvC
vD5OtdXR8GzGFNFDydF256XtA5Kqmh3i/FJzvCD4os1HkcxUUZFolpY1MsdUFsX2o3jFUte3ws1S
eivD02eqayXuX0Om2PVO/EkIPAsGu7n71gH+vSFxYYsxor9cLxG21g+VW9WNi9619RzqalY3Nt4K
qZmqY2f56FWeD1CWkSE7k5Jsx8UNnwSzqP9BGpx+CncjBOqrJtLYWVD46tq7qYNnZLzTLFPufKLg
PLdYRIBiNTprdDcUT/kQht+fVGzNjVpWGTVZe7UrKS5/iSpOL0XPkz6Zhj3y4Co42daPVV5YeJbk
BuJkLjNY1mjgAf7hMjSuowcUIAXv56fYh/CIsXeZMa7rm5WO3A1k6VosDcPfJ/Mxd5xftrmHT2T/
0u35zloUy0FrW5Wvx/EJQHsdscYltNxEiLuHRU22SJWtq0HcEE+ElVZcCv5yndoc5dgsezsPCMZ5
q412CsL9izg8CTTuWHWUCkJRMpfna7SjjqAsZNqa0qn/+AN9myXmLKrRtfxXjweczG9M8Z7sri9w
2uXZ7CkiMlMNEtrpftg/3armEuqfopZu1ujSCrTQIapYk3Xiq0sE1iqFDlV1lb1MDPpHwmAwFMGj
bigihyQbIba7zECgq1dpBXNf24uZiJenlRFqKquh5axoLQ8FK880E03Rfo9yra4H4tl4N0UkazYW
88ZjlrIXcfaGC2FykA+RBc1r2nzUZ69B38TZXg8mnWFb7s5C0LXKMXMNohIkHpFPF/xguFe1z93b
Aa8TZ/3oijMGZXxlc4NY3iUOvtG46cyjAIwyyYx7gOluJqESe/qP3zDwIp/cH2i86NZvzRKSxqvR
PiAwhcHgGJ5TxVB/pcJC/l4tDVp8SRf+lq7+WO9UbqaBpKgvf6GwzdLyY7+2Iqfeq0Sq4D0lkpak
14u9nVl0IEhjVwIR+A5X/QdFFVhypdWz6TJCV5MJvp5qntldihh1/MybH5GC4X1Ray0GvzbHtPE6
QgYFbk5xW90EbxbjKjYODwYKkYSZyJnS8NVq07cyO+ArofKzNyTVpWIndtqeOsTKnF1aiiIhWFFW
FBiL0QOwdDMDNN4YiLXSjp/qrK92VHupwybFcB53cajDWIOt5b8ZQXRAq61osOQm/dOOoNER5Qto
a19t8v/c4oUbN6LJ8nl7XoC0ZqSRX6HDAtUUo7+mCo97RHfaOF/2pEm9EAf3aMZ7OoN17v02sOrB
V13/vjs7MgzuAKLHZWQBqROqUHo2Ugc77dQmZANQ98gD4qW6FT3pdxyexQ8x2/Zbt1kxVC//tcoQ
djyTDVeAP/A/hznZahQr7o7uw324qThyMKxrMtHyHz2CzVm9Nl8Ae37QjWDvLKQ7mjnCgmeQo95j
9QWBcBB/TkDE2wffDL4IJ7boQ5c4gASzSmSzdARtgHSpmQIEfO5Bmn4VceVWz916m/e16VnjrXbI
ANSw4EsHk105o0KuEkcayBjvPY8HDtMTNzHp7eGLHwq5Pir0tlsCcGec3Ge9/c4Q5pbxTG9KDBJk
5CcqUQIwirnEIaXHhF8Brg+TiQ8N74y46766IZkMV8CrS8wFXjikBIkmo9FJxjD2MvVVk1Sd+vxe
vv4M86YO5M7EK9y2l8duqlstwUQIgnk3cMTQz/O2+S5UEtSy0Q7uWzF8TFSzA8a00C9lEBkNSEq0
KXUibaXw9zzAWq9nk1C7GoXmT2N4RCc1aFISj0I1E7+sym2Mr8S8kOkeF5pWtVo25tqxhqUnGR4a
Vd8vF5MJdwJkPTuZP1WKCBbuQcl7QX9fpMWz7ob/3ycdN5FBHXzIINOERhfMKEYCimWKjeHm5e9+
Dk1kxMXr/Fp0iXUfzbKEITvGjVZT/TIC559GAJPjYaOFQ0TvZA2ZpiQgSamaXxRihbOZ1XD3NAwj
9m/6gsnt48VgKKwnEgQBrTqJDpm98d58EQlwtbF3gkQmTArZuqsvgtvNVHAtqfufHb1M1IFykQ9f
71FOdO48XFiClhmwtfG14KXfLYHPrxf32Jcl0vvTjeJvdIMOAM7vKyBk5Y9jBl+hG4zXkYy/0H7Q
ZVj+RWrsLxF9LK3fnzfZ5RrLnvsbqu8BvFocRFB9673fg+T35nw49XMkqdY0xe8ARYMeBD70FAHi
5qsyPc5B2GnNJpSdKcN04KTQuu90sHDjTbC1g14/Ukw2wv9VK8ov1SRWbdLZyxhau7qSdk80tWjB
FKQcyQqniormWo0KymHXCm4+pK4GKgb6bLW2Zxllknsj0YBhF5iN2FRA+mfAOLNEFEEQrHMB8X0j
T8bNT9JMypj9o1NNQ7cofVlxHZUjxTSAv2w9MO3z7BGFSTpGLmj6TwAoyR6PSAV/FmFREXHP59nd
gf2m8ZlhHNIXePxFhkBggaHo5z25ljCtQZJAhoAYguOcYLowk3GfwKPUJgWlYyVytXodfqmE2HTo
V/fWOjLn6lu2T0z2IvSXPtZZwbOonWfWilXXCuatQE2RcihIVRQTo6MFhQI0vdAU6dlsp/VtJWlg
CLpPYBo7oyo/T+cUH4h3S9pps4Azf19TfE7sOaZBON/Hr2mAM7ALepTSgTjXHxcuG2tjyVvhB31K
A5oZ/gkv+VENGyDc0JS5AiYLB6kKYDfNwVhhJDDdl4TyEVDW72I5c0qxEoCn5ogJso67q9zWsYi1
nZdvhHEC6GX1nRWrcxuThVMWCIAVw3rPPY6EOq2Bji4qH+F8R+WEAOn9OGEThthu2VU+2Uuq+RUl
c6ePc7P7/CYDUtVpkcB55EmhnP3hnyakSJoJsOJxwVSptclW2jTWxbKAZf1Q7b8zJoYmWRZFWQwe
CfXBMrfVXwjpgoi237q2ZIBprXWEmsQHoJXKyIkvmzxUS7U18i6v90GU9qY+4RcPkzNeBRp/wixo
rkANXSYBQLKx2TqnohgOCtasvSMbsPwM7wsnGiTWd536xnn2l1h1P2iYBxRJx+xFxJQYrpe9Hknt
z4S3M4FLQzDi52BS+gJ2agRnC00CVJA/cCMpCkN99RIzPQ2CoFfNgQ4CzMDogc3Fm60KjQP8gAt2
Mu1NgCULulroXEA0JxozkAI+54BC6VOArx/FTgQhTy+98RAKwSSowoBPI94h/zbA3ScYaUWIvVQN
23TGcNRVLVOK/VQbs1t8QaKqgi3AEq/ewYRthybcbgerS8ZffGInPYns6fzSWEwaRGudedQHZ761
W7ylit65KPM4xLPegR1x/JCZbFSc3RQ3xpxil4fIEUlYKbNFTxvagaQ+yFkvgrA2kX8RDRh4a91m
HIlrJTujy1M/XIFMfBhNxKPo9A4dtQjbsbJFvoJOyt18Y70bxn9fnX8MN5dJ0vYbCab73/kPOMjj
3als1tJjoFAVcq4g8YMYBnjlt0DOKqlPblsRJHR5QoL3dwWKLf6SA3LV7vAwPc9FcgE8OmVQykNb
lXiqcxQLxKR0tno7kUd0FNWX/kgbIWfu6eY7GU4qipWYZrPTkp/Ns++KH5bvrVSNcn+wsieKBWYf
ZbYgx1fC8Y1n2MhK/KbGXFUjOPs0xUHfCNiyp6Zsy5Ezbg/Yd0+86IaUmCH6NwWxdsUVRbrAEO7b
Qn+ZMC6kIIE+liRkzFYydBoL6aQOeC2cAk98CcgEKT8TnQQzsFu5LUPypx1BIyuIL8UKccStX/La
rHczFf8VuFoJMnjdT6UBg9EOxIHQSdCyGZBYKFnjipI6TMKWjDE15KGFSkSCWBeAEt4aIfS6GPlt
rLJmlBp5G4TRzUB+KBPEUMIXS+4HPNqJq1CzHcLpcVuhF2UQgCxFd0ThH9QfHPkvVY/v2/Wzol+T
iIbudD7vBx0WbRm+T+mHmMNEqrpqIdcPP368StxcYpdeLpbmwrLVphb6m7zqRyIETXtcfL/Karvh
YtQQA+Dl8ftKsTS69JwsitFWW33WUPPaKJxkNR4y4NqhynkmiSpIx3duWhvcqRym2fvv+PlINC4v
hABIIYhHvFA5i09Jqm10rJBEnkF/x79OiYdHnFBpi2PcvnWmrhLcdEqp5oxsHtWmmVj4KpicnNWx
Y+MPIW1HlQ+ft4uTOcRCuHv96uA5rto57TnOJbt4AMyZ/+kupUY1brlrZnCNi7NFcS6c4qJSfqS/
r7EuVXDEDlHRjVSNEbXO731YM9OiO2Ahe8DP/z8I3jfdd8r7uXItOTMQ/sqT/DKErv2scgeTqyGC
22FvHjSeK7KT8bPKVIpUngRRuMICjDuKqQOLAMUz4lIELYbldLLDvJ/Q89uhyVekvDe2/+Cz0k+z
+Jbm0K5vdXToQrpjgWo1AYALN8g3UuU2qBnnIbVE9P+9K3Hi1TCf152JnIb4NZA2vL5Gf3gho6fP
NrIPv4Latb36QxEVvQnjKYYWEqmCzqWazHZ7tQjj72VEOoKXShAUlquruQuUFrK7SUZ/X0GJd4y2
VJyGaj1xosFq2mIscH8sordkbEUyBAgimW7i4a8jx+cbg3IncKJRFUlmtxgx5KH6Gd52dA/Gp5jw
zjezlfeJXMATKhTHVc9tgqJk11bXxEnWGZ5HQgBgn4Dz1oAAZRWQfKkfHXwaf6ZL7Rs5M0PaO9Sk
cL1oAVe6QzKLxrFOqDApr1a96U1n4QaZeQZOe14P3QZJSWRdied3LFzW0wetzF79o4XE2u2Nuy9t
nTLphJLqF7r48xNQ555/bdMO/79guDkcgKkNcWvzKPxvChEsoWq8NwpBruwkl1uew3W2UlHLcsYy
U5QOffNbwo3vb1s/Zy1ISuAedD2oqst0nLCJgSyv1ISSg4V5oLt7Tv98+Y5m9y2dhcnb4Lml9KNJ
12IVAbqpK9d269KeIENDB6aGZ6s39Tjh/JxmnUyo2ibg2646lSHZfdGw3Vw427ofrQa45rGoTBzz
5HdfoKf49CMii4ev5fUSsrsFRYr0HmlXuCMuhb9c3XlHVJUdDN/rYYWTSGX+uVXRRm5Qjj9oFQQM
qJjozDSwPECZYdP8PxjggeSMkP/s5W9I1vj+oTo33jIuxE8wh5xWyj3XmpQmI6L3pmEzrPadUNZE
VS6YiADRQgqZCmxoq7Kin2EG+r8O+b0QvrGkYCGFMXDOLjxRdqkHocxqO1ukGA9eI/R/OIkciiWM
bMCAlMccU8c/Fg8xNhIJqLRmuunemCXB1P71uI5NBfMFC1Tj1JWbNo1bhBRXQ2t/lsz0S80TaACb
x6XOCNLK35+hLp5UmbaN3/Kd4aHuANBt6OWLZHXhL2J6zyCGrtYTwuSru8Rmt6ilSm7H+ksefqAe
3k0iT5TtKaDFYUwRLxzEVc6U6OM+LThSaU3T66j57wVOU5X82GKnHNGTnrAVM4VhVinCU6M0gVrp
FIzCakwKCs3yw7l4xAXA/w8HcdEFvGZZuEoqZylGWKdwp4gLntQSY2wS9c251iDcL/Q/vUppNyCF
q8AUeaz7ZrsZtrR7tpqzE6/AESpg4mSBgEUKhNOAxRh/f3nWJMYg5z/CWzyhlKVM/dgwp3CDYxz0
dkGTFfE0+UcS47ZKcL5q4njc7j8CONszG2NDVDiENqXh/jAEZDXeVK/RWsd8EyKtu6YRvLSbE+Yx
MrllH8ybo+uV3PC9uF1su7WusFiM1s9L98HLnBGePQ3cCnxL0ldmRkMpjeBtjDrKKCarGcSF3K/D
crZ7Zozp2iq9iF7zNDQELFnq05Pu5j+uisBdnRviEQYP6jTNLK/TeFqjkmwd9i6NC/xvAhivjCZS
Qr2ZCaTFIfVoSM5trmL7ld/bDpPw1l4XRHgH7dAni5OlEQ9apMu8DcD30Rg6I9lXYDLlMG2Ob2rv
gx7/BQuLSjQcX6ycW0YoWSxLrmGt4zMOjkncOBi3XjiW9nZmFYgJ/Rivi9wtiljQRIrWIfgw7trc
xKXWs6XX6I3RvnGD71ZwiRqKh61LfWgVfh1D3uxAQa4fLRFM0HUWWjaAQJMILAaJlvY7x/WKvMT4
Xm/umaZZ4ChvxbduQ+BNOtEDe0xrbS1pSuC0SAyTqM6LC+td8N+pY0A1zqbUNTFDyWu6YYpLMmfq
0LqcYVx7TwNENzIgoXWt5gdN4xlRdMGwfqc4Z5Exntc3tCFRF1fxuo7f3u0xznPdK90fdevydDZp
gnPoGD5zLFNNpDwAln7cSDQaNhukwbMAYTFpAuGHVhHJqjmEdlr68fun30vAi07GQrExalaCRyVl
l9IKADYFdI2EqCn7KitlUyD9IQNbi5s67cdeqLYsVcc1JkGKKGSz3WLED+JVqwnYqx4WE5Hb01RW
a/L1u5ftkkWEXtaAEXXny/MZkY2qYpL6cYMFopA2mWIpPirik/Mn6pvMNNQhKNcv+jtQAsKyd2u6
+wPVG5Zv/qrvZ7KxvkYj/7HIDOLKwNOD9LfHDlNDrcSE8hvn8Uacm6hnKjELPFlPccp2L+CrlXdb
Bq8d0hO1pG+5E1zbzU1kPuO7vcSuigju+I8EQPIS/GOOGH+AL/RxXaqOAPqQXRo2ZLZLCOiyxZl0
d8AuY9euaBg5LyC4LXcU2IDzgtpnTyKTEx/Ef7a4U4/eweNzcOC54RfaBFy5izk39oxmdH2PkYex
3z4lq/3wHocjI2gyq+wJoqNTtUldUKIlX9vobcK0Z1yvxDJaXdLvdw3OwOi0RcgL4TjpODVw9YvB
0KF4NzMOSeOR0jYn5Bw5OZ+KOdo5f9yPtQbHlAsDxBRqgGnN4wK5zYzzlQVnHWp6/6/GVlFG6hC8
DuwtCee7/RNRL2cihagbndJvJCAPakwiroBfl+bXNUOUawK0T8yHXOcXxoBMzbUGM+BTywl9l9Sf
lO9EH0zpv51Be0NA6TW3y8KfScomV2+2leErFUrXEkcj4pb1R1G4PMMUsAd3FRBrOqjskuDVGzYH
fM2VTLNN9wffGCsDdJ63BOOrjGzNynKATqUWhb3Ah4MXWEM0QdjACHR6yL43KAlJ8yrP+QC3GwyT
D15/q6p4ToiGU36oLYObkDPetRedYH/zNZN6JPbFfF+5+CZepcXAtXos0e1e4Jpl0hmrc5XCdVWf
4hWSXyqzLX60MqHq34a42z8B1C9LcK0YH6heCNm4bGrAdQ9Lr4GlgIAyW7Y+oII1CMfmR1lBajHC
JV80/hppuHitE19KW93GbafLjEgNqVi8cpMn8OgFl5qbELRwHn5r/GIUTvhhA1q/V/zYEVPSoKQW
gb8kxJUurZ4wgO623FK3u1BpZ13B53HReojBgn0TvKeM7ULSZxjdOYhz2C0XUugPH8/v0G1fcNO2
jfLfDsTeXMFEuamCvimkfxHz1JkBuxP31YAtrIFvvYCziXbXdH1ctPQpGKu1oyB3xou/4TaQgjLf
tAGdyadMnen3b4j4SHfA+hP9w6KxWng20Hd+eirmF1S76QxASxmCN/W0zaIIwuiXLZUdiAFIPX54
f0Z+uxyZVexfYAF/TDpHN5HMripAFfb2xjdpgD1Mk3yvsZ4BaXYmVOYi4opQCoFTbCwCMw+rZ1Zm
Pc0zLx5Wna6JVTxz0aLuQIx/E0+OeG76/VKHWB+POD8Kjngl9lwM/hUmlO/CFwq9s8XUNy7iEsja
081F74TaBMQYEG9N5XjI8ZbKkgxrI/Ci35TROA8pbDCgDFPZUPl2VBn0YY6rJO36+eO/vKQYxYDS
KVIDIsko+T1QbPdX58YgwBHMG6j2rHAMlFHybmD0uZajhHH529h0qUQ8IYWB7V+NX84yJ5jCw8Pt
g9NzidMinOxQFkxg/gfDecG9DyctZohhDa1pDpy8rvigZ+CbYugPSy3PShelyABfYPl1h0mEEkd0
11/G7OeSoG8ap89DjNjrLc/DWgREKqbUH+a9KWT59iKZaMselKaD0j0X04HhSTHdd+0IE6RDfoov
lLSRQb3r+0aBtbkSBnvoLAkR3KRr/EmOvGg7rpcPMe9iY7GIjswoHqzVA9jLYH+g2ODysl+l4gWA
mWcTw0klFMjEeAVisre8YhsSG1qmuLKLyFsJzYtchaXwUYBVtJzY+gVO2Y+zCb3SQXsQu30Y5rH3
5dm1gJhZ1cW5XVANXYF4Cfe/GkOw20QM7M4pskYf7eWmv9hOp9I4QRZkT6LkMgXtL3tmoN1Ltdlr
ssWAHAQSKTn65jmzD2XRT+QIanDJv/87CTkzXs3hrQpvLkJF3H4WUeSPyEcmbzziOwgkw/a+Z+In
AwF+Gc1u9/yQLzCZPTcs+tzCC4JumKdn2AarhCiKlAd86/QDcR7cfvUQuB1vF8MuM0FBnWeYyAGA
A72j9yms0SgFDNSD8dQlp3Jf1jZc8MjfbjxhWDFleHbMN8A7RtLYeSTlcRd4tf6pcrfMdnsgC5r3
0lXCsVPnjYbdrJUUX9uf3pOGk0FJK3lPymMqnuNwH2+Zi2gEKyRRjOhpC7kIc0ylt6HAEEs6oUFa
LDT61ALMvgiYiDKS3PVOf3DaSnOdQB4cki7p/JtvJMF7KcvCcs3Id0JArRpjucsm0xp12nhSQgRR
hRIB255oRUqWys3tGXqlGpKykTll+orb1jfX7lgyvMJZ/Oe/hY5CJ0iyrWHGV/flXR2JSFo4IQe7
AKWQzX6nhJFe7dRJv1KckxQN7Dy+oCz08xle+y6gvh/zQUkHv9UVy+y+79a2eWFDItWAf4As8br0
idTMYwM1msTliNgCc/KP5zHLP6r/tjoakaiUb13gKAdsbijj3PVrBjTpD0xLeEUjmpnshn5g8k6a
vo2wdb6YiY0dt917KT4pSLf5EX55rLFPXfgXxOFOy/sJK6pWMGfjCsm7F0t7+65XM3bvgrGEtkjW
DZQSlZzVeElPwIEnxMXnRMTw8dBbvkGUSaelUw3IPEyCpDjd0aKhVIRI1RlhZVJk4s6JnvnejFC6
nwsQ+2nXeRgF+J8w2MaG7owxYE4923BWHbxdCTJCaqADRyQ6DC1FU0YYimUvryrG0649hWIOvhNq
TBMDO6QSOe9Hz06kYiOcri2ZSBFV9ZnnhmnjT1Ojge+LHcDhTqwFLwpGSX1MujhQ0hL8iJ4Qb7mU
eD6O/cYB6Thu0SyBl8ooLmAHSYrZ1j69fqI+q/u0DO5kM7JK50oH6ex6nzv0Wlcxy9QVrVGrCx/x
5oiveoyvNr8vsngbCL5gACAxXTqY6nm9qEuaBZALsH2cJJdFNcOBmN4OfLM0lNLOUT9UhnxzJ4Yu
B+t0pb4ZBkVQWa8lsTHH+OAeiov/Z9G1HKEYAQEAVhT/9i76S/fp45wk8WhNoP2C02NEPTez90Jm
d4jfuvcNmgtHfv2g6hqxz2M4XNdIHzC4SxdhICym7Y63J8T/l5pu0wvH4a/LL34PyJJIWDYXLFUW
+1rvU73d0rSa1vGMKKTrN30z150VA5PuDWycCXUTvNyjLGkEQbvqaebmbLcCJxfhytIuEh1UipEQ
AX1HK091Zun8yXZe3RKo+3cd2M7AKzh99O1ALKgr9meQ2absaju6dlcvTEulGlvHjo0lQdj8zGR4
MnDOMX1NFORJczicXZN3eF7CUUWdu/SyFz14DUJDFqFVLKWCaShJXNb8DAFnkNQJE+m/PtckF6OG
1y7HvGLV2PRIPCN/Sk4dbdZKsct4JoIh1oyUKPe10ro6mqEW+BfVxguSiIAXs5639rvTRWw3nkNX
+yS+jdj1VHd+8ALPdivAwJuzF6gOJJ0SLZ2GEwIcVFoOkyZK0G4xO3+wK7iUWvUljHHAzGbN9BRN
0m/7lbwVNYHx6TaDR+Zcwy2Y6B09XzPiajKk6XCmOG0iAGSN9mEHfnTeQm/6b0Vv+3dE4kNbD+Ep
afLRAG+xNIZsXudj0vh/arkzcr2AI45/5UxJ8ENe+G692bdLOgeM5iq4IfqjXK95HPKY855pKH7V
8fqhz3pBUFO547Zl7tiC9jpupFJqz5d9lrBG0xcsBT38lo/1vdkxKiy4tHeoA81ha7LTjXu0M+yi
PMmZjretF3KsM7zDhYtIFhRC7zFs5LNzuy4Whqjpu0CDYatVuiftFdK9NaeuarhXGv8/Lf8w2szd
It/7Jve4jMti1r4LxPp2hdBbzPnVk5I4g2Z6VWpVfB5ALDS8diPsuOorM79XQECPKXu4QNQZLiEJ
fCd75BFp1vEvOBDJ89szQYmJlZmZZlOGzD64P0TO/Zz7xWaybaNi8PkDwrYeDDQ5bWENW7Ma7nxT
OJ6orpVncSAJwuthMsRCvxrG2PPkl7dYyTvEDaS50TntMfxMQaFZv7Tf8HK7Xe5UqG4mN0LKdvtI
bJo68qaNWVTWoUTr2V95FvCnOoucBDR2K92pcuFKnqy/7/Ydl/OjQj2BLCO0mzPe2tWe1l9tvIoZ
ZCKT+INyydBQMl/+nREmW/VnSHc8rc74by5bFNvAGKWZE/Otww6tXBCbF3HboJqttO6luH7tEQkr
+GPG6Gk6vob+TNTLp3is43aHKvDI5z2lv852k8hrUNPmJlBuPH55iMDlR/xm+a2wXwF6RRJwG2YE
FM6m49+AL4kzsXg7w2C4slXDiX2ms4eFstRq7bh7D6GKr/c9y7rEenWiAoGxXyY0Xc4pLC7WPipc
C7U1dOjtux5gXzzGuv44g4Nm43EXbxSd7liiCtLfBO1OZP++xICYaC2qlQAh2c4ifWhV+S0iOIQs
Mj5VjVPpPGIekhtgwIDjtoxuxPrkaR4sSeWPfPOilijD77eESJHuvYyNermW25/I8WvI3V1AH9Pn
9iXLLv7CcTxlvCZn9lDC3yGBMwVgE4w0M3vEH0GN99q2ixCio+HaKp6rD15sx+/tNiDuSfZXbzH7
pOpq4wzsHLjRqQNXhho6R6mMw7R68BDF9ivHYTFjpFukS9aaEQ6scN5hON6S/1wxCxaV54cM6vCG
hrKS2Ce9nHLhoFScp5EkVkZkjP/0Iyfo1fSwOCYWwpjm7RItsAGpRkhUZEbBVJv+TanTFu0oTEUv
8QBPoRKAj4XD2e/PyqKuNVdfqSxFNdYQut/J297+UxzJWCXzi46TKgaBpCWnr+z7dgM9Cz7D4krc
vsDFOVzgF/F6y4MLYXsc3/6SVz9YXQKCZkhf8CTb1BFFJ3TNGVg2cKzjpsaqiVhys2vDSAgBhU2Q
p2j1XrnIUmMq3F67K2+OE94hJqWJNZn9wBpwsVy/xGAziZAJrNExzKtxNV0Et5CTymmx6evwsAek
x/DDYEA7HU2gNpfwma9U5u3W7zrBK9R+1+xYfnUCqAfYIOXPPuGibKFtPKB11k2mT3J7aLw1o1l9
WKBHJgJOZBxw+RoLZXKEW1srKgGrgw1VwMowsUJy7oaZ3HYczHDXZ/f1D2uTMXonmnxB9ZJ+K/Wr
9Q82EoQ5IfyClZhmC3wnAqepydyKH7HoYSYwGjLt9FDmTRrMuyeXYxFveQpuBVCPctPQWpf9SK0q
gShdD0C4YxS2i/6B06EctTWYg8c4JKx48D19cnDqBP1/cJ3EY2uUY+GAaE5zstxqT0dFfGef+P8Z
43b6s5cc/yONnZCPZ7Us5L68RBeMYWws/+tmWMOwvXMchWhcc+FxVw8oQAxTFCjXC6bxHxp/RTVA
VPKUH+sckW4mnuZHt7KjgHyDSi/13fL5naRqY6kRsXW8uecK7RB+TvmFzr8DeGQhmOJBPfhuC02+
lNQ/CfsGhKsC9eRSFC7vBBGIdA6jmiiQ90F+sS5iR2GGIhEKIXgBTyaZNVW1gwdj8o4lTMh8q3pc
fn6gug8o1S7gHyWfeWmF85RLcoxXsCWjpEEUpDPGc06P/LAoTw3rSsrCcnaTr0KUk578RRvko5aH
tA0OyWeDyvvaI9m3BqFajwQdMOIpvhPMw7SJqF0i7rdhl2VpF00FyVbd08u8zSXcK06+bZI7bP7d
0oAOqfZ8nIDn462LovukDIxf74Y2nPCNHOJInF6wQLUJBUHs7gAQjvCc0d0Zf8T26KhUnMoQHHnh
NMrbEv3GVTLeZM9yZdN7FxVeClIk1ypsywaDV0UkpVMdaVL9FSf9w4fTlYJqWFbYeFT/ekfu2ZAA
qiLmrO+cRD2JHDXB1SITdsTfPyWaDzwcPtI3ECVVbCNkFnwpKnoddDBvonN0JQLrQ8ghuahlwg7d
P1xeMT6Rcl7eDlXzJxo9znnlN7ZYCqVml7Mxq2IMaB0+vEpLKf38anivD/DkpLrwUP6JCAhwt243
FBUJmbP2xCXm0YRO8Mfj43ISmAnDQ36TqegSbSYq3iT/XmHJRV0Al64I5vollccx2N3hUCe6UV6K
ixfMo4Lyn2mmNoKiwy2pj+ni1p7mQspbpFNzK7JVXXUZ8WiJIiCyGwsIbuclWjjiHfleqTJJuLG1
EEj6qmeG426aQYZUBVAcwbGh3a/Un24IHsQ9gFOxdg0gfCRYZR/GTtHpgBf1oiwmYJ+8g2OaK9pY
m/27YHmuYk7DBCthq9pCreouCBD7bROIPw58AUzw3Qa9gu/RhlNzoA/WN1Nw7CiriyGc53LOzWR4
0w5e2t75vjy+0J3IxBaDI4JztSL2rIWGZfluP8imSOl/i9VT24t7FBUTwrlgo6HqIHu9x0df8xhb
8AiNdxUa1xoxSrbdF9zxp3p8P/6LwrqFVhmwCiEuzmu19KPW4Gy2tUil82qg7VWeXl9h1C6W+PHT
n/SjlbEgvR3rMNDKTDPtIEDZpntgduzBlyv5uMZPQrf53y5WP4R/TtXYqCGBez+F687dkpicfnHz
bPwjjYsDUWyvr4uobYPMFsQWHDhTKO+59LspBk3tQ7lomjUKKlzlfnmCqOZ06eutPzTelXl9RyGf
FqSUisWQwdrzD5Kwq/n4QHGyrH4HNIgTDI+k8Hb5MjwiPmNi6/vyI6H8iKAG8ReCav8F0i16vM3D
ooIWWAbttqdoLIHJsusjT4d49aatmFdWggTrOSRyz+yyv9fOPEZ0X8BNjD5yEqarleM2/ztK9QSr
Cs5/FSrAl1TE3kT3WNPCle6Nccf++cZLOyYcVqfAakZKo85ZaYyNfuq2UnDUm5bstuMFsq+voeVo
0TJ9ADe3nLzDVT+x2vgEbCnO5tSQn7JyihuzozAcNwj0e5E7RUGCOng3Df59wYyYz0VBZvQ3sTtU
xrnAgNqS9vrWhmz6ee6sjNr3wFjoY7e0THtxAQcFdkiJ0P8R1KjkmpO2jdD/9vWj+KR1nk5goFfG
HlMfkoj1knNi93Mto6lo6/zxzxXqOlwA+8biyP2Lq9+4QcVZJkb6YFSzj0n0CvSPYTLXJY1vjPDp
Z+hujp2H5kp97mWyNG/CTwCFevEsQf60ojVg8r3dXtQ8X5+qbzOk4UaE8xWJPuL7XFhqWgz+Su1O
DvopSnSLSWw/YHy8aa40m9WsokYdkkMWBlHVW6RQlKvSGSPk0uM6xKFCkQRYLkoYTtaidtJ7x26C
p5eXgXOy/V+/CyGy626x0UmGF7Io3xjXPqP6VC1n+lc/NyFtIJpXyjOWA87MhPR/NEBCdjyrA9UW
uy7zLFoC1sEE52VRKcOHSA/tCE/2aEvylYgswSNIKo71AkXuytPtoujhnJ0TDTxblHi2DZxf6Ia2
wM98Y/Hh0dcWMRO6Vlz6XKTrtmkbHkM9Lw7Zdeq5bu6iFP5RsaehKqdJ6LoUPOhCMMyPCmF7heKG
1x1Anid77yqKCtrcNZtGl2/sAfLKrEYWkcQp7UqPWzYo4/fgnF8rZOu/Xx5WaVrRHVA2i8MTmqjo
QnaIbUFTMkwfLbDlyoSYvfmEk9NHbQ4YYWNmFSVQKdb5l1cpL7F69d68B7QyGfj4/bspe2fv8tTi
NhlqeDh8cUJ2IpRiVC9Z9AYF5ViswZg1Sn60Vqp+fdcyw56Ul+ZSMiEuEHiGr7CaAv8Ej61Kv9En
qBp2icpD3CvyosQLS2ZFN+iIjZ2sc5QathsIj+Ofq9o55U0qx7MQzlILWwiGaE/6dKVQiNrrPrEZ
B5XxPe56JCJzfUSORjfrKjOWfnKbL+8v4iWPlYicahgvGZAQ3j/3YtbgFvVECEpLSWj3DoZ7VFQe
OvD+wJXBN2P07OaXPVCT4uoxH/Y0Y6Fsqcxc6UzWxY1SnYF+bU9PCassrnrhvzV+WL9mkyLzrHWZ
oury+SsgmF+2ry5YaZay9WhATUdQ06YhATzTatt0p1RaoeUG7JpdGdinPf4okIZWgPSqpHMbSdqh
TnxOp2wbTxb7TqfcSgZL6o5wjNcpflV/r51NVXewi1/kjG7nUMFVu70UbP95B/EHjnI3WA6viPOX
A95e/wLIPSUQLAZqvjenKWP71cxS5apud1gLeczNH0Pz2BvGJSsga1j52J4xeQJM3jUoJ0NBBf0o
fGkgk4l5b1Q0C5ADXbFa1yVSLtdH6h5+VRgliIzuZvVPJjps842nNpIqADNNXeLwob124szwfvvm
BpmhRhDhq9zGWcUbJ/D65dGiHVe1DhN032sb4yID88MJqCKj1uS5PlkMU03TAZY0ZNshMWMxecNw
Zz9WEG2NJRmtQ4g5PMe4H/2ABEVbmunA+K11VyqY/+Rm+MpHY0nCOdCoYkFRjClc8heJPzzB/N7g
NEewqcaediiCiroc4/d3jjyggX3N3CkQ9ufPh5fwVsbzmb1dshBJiZMFgxLBZWtVrqOlHxiuPcbI
/0zAfDkJiubZQw55U85tlFysZy/wGS8utVSHDww3rltsELtJLby77QXMWLcnjNveOIYyR1dIyxf0
V8DPD8yDyMl8dI74/2EKDpQnRzQiK1dpapvUTXt9w/zIT48Z4QWnIZUPNdCe3nHXXixmfp6gz/cj
b+QiUwB1uYgMApo/lbs6bS8dA8MF7pnoqJBZAQT0A5NT2sL4SaZtPIYFovtSwzyxs0hgS5fGtsb1
ia1jJWe2WlXgEOTanTPTxkevfVWGziCaAdP3JpexcD7RjF7aw+4r3mmiEXd+QGAa+7Yf5q+k2/qf
rHB8rvkX+V+yuLCJ11Qx2T5KkeHdeWWnVFvM0x75gkKZigX30UpQzipGTHzjFV/jWlmfXA6BFLhF
FXDFf7BspKDjkb7J3H9Icz9fg8SbA0Kf/dJjVhGecQbfNbwYZsb7GOLhgFEbhWdipq8riG8D6u6p
H2rXdvkjkeN7v3ZO9O8oXbJnPTzjpqgccFFMYYIOhNaAioFvv8CVRe967MvduPTlOm+jpMPUM9fR
/lIIrYeDAgjN3hMSmd8tSzn+cQFc5l2J2gUjlGL8mm/A3Y0uA72/y60ya5+AY5dUEwbFZxZruFJl
C7YcA5o/rGX62T9nmAXeMjgXzPET1pMRK/IpK2nfBrB4NI3XkjaIWAcYnb0BwR3AbtDk3eurCEhR
KdzsO8yLncv5zjlLO8pSeT1jlQ1Pdbi7yckfmRUN1Y3dviv5YK7JShTFxPEowK2EB4opfGcZfYDN
SVRBpc3u9FzYlOeUE3oHYqXMo1tqPUJkXUZkNO/QmSOgCr1W1kRRcTTo8VN+kOKGgJfyyQ1XY2/w
q5Aq6WI7Buo6+nmPGNntDpKhCboxNxcFP3ML5fs/GSTZDOdLr60XcdSswNIk/Q8+9CL8NC6W21wH
W1oKavp+9TC0tVp4xk4sL4wYvbYkLNL/UdPaAFiSkjzSrtJGn+zxFgh0xptu4Ye7+RG+9atCEuzk
2y81tYDMYyyjTIvZvH6pwg0477WAvqNGzs0/87Ho6HwU7uCcrKqFzGpCR/yvMFU8puGiEFNpwBTE
pem0H6rKB8Dt5f5Et7oj2WnHnPIt6XfD3DSFXA4/wke1cVACBWN5hDNiz/BVQz57ZgV6HI/xB+uG
Vy7UPSTJ4+afrHSlAJn+D5dhm2J0BqGj9qnZsMkvn1AX6OuVYjcd9LzevkAmLFzjj19fHNUrdDTn
0XEPEvrwqGNIjng+T3DbfISaNZIWSVpzsZ0e38rGLHAzvG7n62NAPbvUYaohS7k5uq80FqDK0Bsb
ilz4tYBUfiE5jFtzz6TqPgn0SelCuIw1KphOKptGF21Xb+S1qKG8EgSunDmNlNxpV5e/k0WlIJC/
Rfw/84bdFvpkCnGpVrEVyHQMPlADzTWaROyTp8ilgyCb1/Xd8JG7VQ07xuxgiXNn9gMpV2vpudvI
Ml0n+49AUDQcwc7zWPNugivtgcYkRvIU8GMBE3SQ3vnZ7pD1pupWKWDfadLzC9Nd8gVDihMTAgEP
gNXaivPAAwpe26MbOzEYaf/RQP+FOsfXbLD1+6/i3HNyj21e2klXfHEcUPv60Ap/N0pLTXqZGg8G
U548O1grig5Uv3sDvxqNMMFLIF/PHYvIdn9qc+sOq1Pxy/TnXfuAra2wvwQ+ZCG5gLdO67EXTmQn
pvdxf0PfqhP+kND1ccbCY88o2UEIlzaWaVMLBdQTGk2IAH+U/SgYZ7sAivUQRa994XQ9gKPqvCKK
8h/C7hmhAvpuHXepbv8+BcOxcA03eFInhRE4E6SHxtN0wFFkgSGtcO4GoDNRec+eqyudc4RwW7ee
EYwwEvTDNh1vfrnphTkG9WvrZ1R07Q0xd56YiRe19qrGVmLWZldECf0tMAMGDqCEo3A6B595AChv
7fVWnVkb2QobPMBpICf5eTFsKe0cvGRLwtlzt097Dn1XO5GKXh7pzOVRJbrKlEnoHP+2uRcfLW5l
PVNCXXj5F2JGfo6dt3hSfE78MsJRS/+xKkdhcZCg8a0BP6EhGi8zLtR0XDA4MSmjjGFFd33cs1vh
icKRmBY9jq/Jdk7objbp9BlMvbcJnd+4yPJ+GATeJQO8qrmr2/2RgKKUdisNYzxBgzEBDXIr5EKL
Nu6y/fupyXfzwi64uNriuOmv1RDxudj+j3jeRkDXOrRlkkNwFSNf8JskDzrnzxZkmeN4yIF5Y2/h
Zvf13qFpvnwRDldW5EzRFixR9bnRpx8cA2vlLI88V9+aGhoOyQdSkJy8iIZp3Qvh5Axm7CBLTsta
7zxvciyMRyguCO0Bc7wjQP5jhGyEkj7nJ/GyJbWC06TSisGzunaKD/REVKxOi2FKqgxg2DEZR1Ko
f3o0DB9AtQVocTlHV86sj/GA0CQ1/GQdeikYH5rzccaRB4N2ApL2H3oKY1ciwRXQxrWyiBP/kxWt
krB5T/lVwpPYjqO8PnPZaVc5Tt3yJfz5qeRarQWle0SRuIP+hbqKZLj/tofRXzK/3X3BljScQhln
KgwdzRCUDKOqs/69T2unqVuHDrM79XoeWHhSeDSRhgdItbPElGPjfaNrwJHT0uA4LD1eMcKVum/h
cyj0nzugjo6/OcMUOvV/LexpVZ9NrZp/yAt5NHXfWgWxV20HwMQmzRJMm5NFv3TyhGlY1J3K5C+C
Qzx1u6xqMuWZQFospYqXCCO0bagxSjSAZ2PeVVJEHQcdYrx01yRwgR7ZQdRgiotYQoISBWtl+Vn+
hNX/jKZ+575lu34z8Ar7CmzeQsP9Hb/DhrzlKK0obbmk5IZfQrkPUUYWuHYRCmJl46F6rppW3yfb
YPKyEDvutIBmpWEuWwYC7BicdKR6T3t1mQ7jHQ3VVw6us3VDHOB10mCPIJWasOFWR8lfus0TePBv
s0ffMCX2++MceZ2ylWr4ukU0+jgDnGvg0rNZPq286Pa65rOkQMb36HSn8Lu93PcqwWCye6Dii4Mv
TRYDIINSLFOs/Yu0lp8Wfi5MNilnYfyZ89UqjI7AmElnaJN6Nfa7OW8c5hjI6EqqIPH2TWBasfxi
zofOHCFYb1x4TtuwjfzbQsF7JqABb5x3xrCVRoi3/snrCAAmXIkHiAr7Jx0/ac4VM+fyLbLxR4ph
fle47HDnTVJJaJmSTdYZKfx28vIwleCVvA6L4wBVr+MwTlUXPRhm9ivD9yIgm7BCmh8YadKshvDu
RhOBlzU5co/a0eyOvaGw/ZaLw7J27N8CvZPu/kc9u13UFVkq6EX40RMsD4CazIA0qMb1yzgY5fhX
rztIHDcjaZIuP/UYJY6tfokldHVnR1KlJ61l8uX3osIvTyDiE69d7ZkdHFtQTUHpN2PIYwBReSQ7
1x5WOar4z2RmvSIQXylj3AeIYncUf1yDLU7xvzTyYYjUZANz202guZR7I9wlaTtzBBVMjXxfJaHB
J3V7TQi3ld8PtqAzA9iZ1ae6pPhKdoq+Sx+gR6yrD4kbn196MqEu5BY9CGXS3W4qq1vJ31nui6Zw
IEdqKZvegDi/NOsHrPnRhFfedklDeWUtTHwn9PpnoojG99Q0CWNj154c1uVR4CHTmG+QJIZq+3Sd
eUJAWS358IFy0DfP8ZPXiyF6NoLRv2sx3qePGbv30UQkbMaXNN81C/oIutKm+Mo2l5sBfcnI9Hb5
cLHk1Vbn5yiCSFYqJIVNyZeJU2DpQeah1Ycqta+enPOFu/g/+vGbiK6xnxi1JZUZ2IgUXQ13odHM
h4kwUAf86auap68NaYVPpbblr0EHkaIz/I0lQyMiXCumUUGjQuy/p9QNZuBqBDnhGzNhJOJaQKfX
kgerBkxZm8RZjv0smFB7TUkdX63p4t4BGm7tPCnN7GbQYQtYtQX3MQEba5Mb/697WeeS3IivEtH0
xXbgXmLTw3KsoYMbC9zO/oase8iz2CRfobQdw39bfBT1+i3sB/qH13HkTkgPIoEYzeK5k9FjXbdu
U6U9pSD+nID5I+qGalXI5tzHo5WUn/VCU2pNCzceQPYtOdJUD87HpVRBPQhMnDp6baNA9gX2ysfJ
kgt8k1/8jIk6W8Hl7gp47ePoVrNJ2vrFIi8VjsGru/XIiF4JorlQImA5g/sdcN6PENwgoJOgl7f5
WgkocRcdCoCF3AeDPOCiUdezLOEkA4yvdyVytypxfhnJ+wYmZLTLrMjv1913BdVX9ZqYbPvKBQg5
Vxpwe3qNRGEBmuXCO5RBPCp1KHwPnkPAmULChUwGKQNEMutV4HVqGl2mvT/zwe+WVoyfdIIfwldV
Lp9JmxoYqfOCNwChMiRV/uTBkiHx3AO6E1+Gn+sDMSliVrvdQ5rlJ/SF52jU/0ncfaunYwIw9NK9
4oySd2h8nmBbAcXc3AOT/ugwVFtlyjU0H9dOYMc2u7xKv8QFXpMcNyc1XTrdr8SnAYcDheHb2G1S
ZLH7LZQhQ6szMB0WZyThzVG4mf3AFa8Og8dbg1t9AuxZli1aYzDt1v5r2ugE1AR0qmJoAqpzCOoq
3Bp7P35f8kdJs87twjbr8avo0ZwNQ2m6l8rZZOcT6nE9ex3bSMfBnmxmFbjJwe4rwJLwH+3YI8fT
VNha8MRNBzlnuTTiiaHaA56uSeKig3TugGca7mamRSB/I49NHcdS5sBbRRpOkV9nqnsG3YyxywQl
eZWnLZ3FzjJjQNvEzWAy0dTF3r8YQPDoEItPfMTjBsBfz0QbKt2XPzppi0+GA0NkeCxCGLtuS0DE
KscNCVATPZO1KHXgk6w8uBz14DjlzAZ76T4M8xiKXO2cIML4iq4wU+qIvennQNdmd92kPGSnldK0
h3rdnjCSljZkBPviEiQ8T8sQYgbRAMWL+7ZUXKodgzklsJ3E0ZKsJ2vyraV3qiim74g/R+RYnt/V
eQYfzLO2iRLMv/+m0G36Bo9AE+apadT5G/NI/gwuHLoQRvGWyh1Vz5DxXAF7S4Wsp+ilktNDB8Yf
uiQb00FYuAD0q9NPD7cxKmPBfhgiLumtRSPL2TQW648CWUHs14Flul/VeCtWDLxUXNzhfLh36whs
ugyWyQpxzgDA7YbMW+TCV2CTAGaVENCx4g4uhCI6+VJJcwdqviNPe15aoNgNswgUgZFfPcNeN10n
5AdWGln8dymLBVlVqKVtuQRvsF2eOY2u92a2HwHSvPEvyMapF+TlxKYfRRvIHtjrlaW4xrAJc0If
AhKdEuJ65Iyeq1Aa09EDG9ZuriTbiPvujUj5xPglqCPwCgBaE7OyX94WgoCZAofRQAH9p/5VrAAQ
q0lXKSEUpXWa9QbPgi+IIEBMwYZOhP7MGZU2tFi6dr2RuW6AG15+uBtypZ2jz08mKQlQyRJTI1zV
rcSw0cDlr0H/xwlSEbyNFnstzztMLACyaLPqLfVLc+jnrfq4eWZumIHnJvuz8E1pass0Fj3iIfn4
KXHWXSzVkD4wvEy98xR1Z0UN89dPx28ICIGVvJoYtNmzff0t1dozeeEWKblwMK2/2moPB8G8xNhC
QWs+9bdP/krwouMi8/1D86WX3R+q+/hF1DSAD52ULluglLCNcADiFHjwsedrZ/fuaccznntRxk2C
sfWKe/o8yBwxRG/QLo07U9IcqLb9itAwqGZWzMfHi9B0QWsQ4W3PUYZm7/fQV9uUrpVLlgTtWq/m
JUPR/+0oPPXGZSdzjEY3e1OrFnd7rJh3vXNnSapppg7wYbR/zql+Fa7Dsnfx0yOD58kC0LL8zQzI
vPn8WErrPqDjHmOi2srinMSHh23OUeR7AQdg5bSkoHjX8yxxFZpJI0aQBYGGAmj2937GkAy8g2QU
GBzzUqZfrrpJ24kfnk/H8C6gb4wRltRkwRB1uWxt5Giy/6kVPGT+AT7LXWCqnHdnVp8nomx+oaye
qYeToFpgRcRP14FAX39u2XVqwajVBC7DlY3GNgrsx4/KDM67FLnKq1Dp3rpJ/8mqCNf9FR1znU6p
oRgUGkZNmlUqTarjH8j/wKnCrPUBKmft1qFmzRR84v+M9argeen0Sln0PDWDU+tvjNWINp2YY1jd
mSxaqPLV39Aoz08sMODoLhC9dRfIRzKUwtik986ks8L04t5KrxiZVpp/EDSL5xJm3tmxg3a950J4
1MsOtW7JneFduxX+/2SJvyvfS6H356Vhf14aiGqptqtR87b1muL5fIAWRHvSDN5CJDVlqk3BbGT2
YH77XMvffccW2KuUp/z6jWZlVYA6vVL6sq/LYQFIEHbDWpW5ahHmEshEsJo94UbNyDfVKA266Z94
FbqSe/1iMXKJNZR7N3id99HJfVfl0kp9H9EcWa8we+wQPxREcX50RL51IM8LLXRD66JhK3n3nnmZ
NE29hdh5YVlZ/Dwt/c999IySYI0wy4Ozc1j6sjMHy0v/riwVQ5GayN09T/xxLAECbXFF2v65iEv9
O1ZeXDctMG4YBAa3OFhNUH25CY7y2nSfN4qTXZ7bZUrpdQFN1H0jpyS+rK1jr55P3g/xhNGk328D
bUVQObQXZU2iLU/cCOZX//TTLtKi7VmaNy7OGKob0Zl3N0MQGfL7B+TM2JZUNh1VazpYBuTbKWDQ
4sfjyBY7aP8YIhTdQOU8MrUVCbD8mqSgtkABuZeU2vzJtKKKEXQY9UasW6EHLrnAXrzSNv6PPHGM
A9XqxmCEVqdhatbi+ycGmTEcky64U3VxIOWTYsLr0h6KpO/h28ZBMX8qgQ0ii3C3QRJcWOMGGKeX
XlkJJeQLRBOiog/4ROW6sZV70OaeHH8S3rlOBMtSEI5hU+dTz/O4yxmqXPXBO1h1gsHBOJJn3XU0
VDn3XFL+Mjb5zoZZ2gKAdhKnPMQ1JGmLG7D54gWXFVH1VcHYgwdgPFxmPWnAmMsqvIm7x4ZRuhcA
/tRKvKxBpm0HF4TzboGUKrGDRavbYxHLTfE405Fm1cO9rKNg3+JpgKwUuIfq0i3kHJSID8czYQon
B7NQ5AgXpuM104L19x50w2Fl3pXog0MVrqjmwWAoMrBrGmV9d1IJ4u1q7C4TpdCJeyrFKV5jG3Na
q+pqfeNAMKVB5+ueC7jWbbMkYAyBiYpVhNXdFIlwrBWoOfmiRgmeigyJEQOMdAlCg7CqBrxRRPjr
kTnTd0VWe72xVmsC6K1fxx9wbGXGmGSKtBWaeWBMSAauH14yuf9xVcDfh5Zt0mpwG1lbnQIo+0iw
egxdp7ablGXhXtLRTsq3hHm3GccFzp87VJhKpsWqg/8PWEKeFzmm8lH6KfOlC32bEzoT3kl/xZ/z
NhqIA7amKjUi998NrS0jUMALm5NwaInTZTiAkGl0HkU0xdG6sMBWS9pKyTJ8uY21/BlYrkEcGrS8
D3EmHAfUCiyclFKYkJOTZhRbUxl5zlQH75rsIw+WBDgyl6zWHqaO3VvPTR9gC8Kyd9WN0CgDJxOJ
duqa6kBn4mHTXkr6a1QmoA9qHdsoJU0NCf4Y1qDvP/or4nFXCX585XSpOX7HuT1X7JpGTc7Urtlk
zFcJsZHwmvoD5ghiOFu6c7dqxoi2z+m9vjj8kD+n7v8KTJTlXDgmvLPPgLOi0qcwsGy1Sp/4Jujv
HNWtxjuQ9XS0yiFXhK0SVM2OBpO3zXJT6Ea6CpPekWwpaPDj42/DZJf5e48J4SbqnUKujoiKJwbj
yvg1Y1FNz8NMTmwnZZuc3USlNUAuWMFvz+hwvo3/Xc090zjJPtEioPAH6l5namZOWJqKABtZ1bn7
Ch7fCRpAI+nBhnT62rnJ7rPFzkupq1Krh7q58sVoRUfgpq56gPRAzXtRv7AJQkY/IZzEutCOZE2r
9nTrQdLHHn56zokaNfpA3Yu8VZx4m1OC33O4ZkALB2ojjg/5IL9VIzD5tl79toBnYIVPPWkecdYT
kNzUn2vfO9HwfxXn+BUjI1eu/IwK1whxRixTDCf20YNn0gcUJent8yuq/L+E9+nm+KuwSI+5Ysr/
l3aGiVPj5FLPG6J4DI5pkBlcopy8rymatqqsDJ3JUM/Jghk/fQWT3dAZMPjJy8WsrYWc4LHkgdBf
cnL1Ye7w7AkgLQyXI1DoJPqS9ChTVoBho1SU9lBRPGOHxOeac1gPmfTvc9Hstan3I1khTWpCbJsq
WR1Z7nLcEfpB1BYScopacWQhwznwKB8D9bHv4KbsILYfH8FR+kJNDaMnD68qxeFeLgQSCmBCEvfE
bNW7nzlceMjECOby1vnCs1dQNpLvdQAtLAX9oy1xRuZW1Qd4zc30nfnphOvzO6KKz/Go4uKAmANF
w06HNnlZd6kOoCTjorodWKj8glWB+SaIT4dbHvGc6h1NiUJ1v6nzZsFMOz7bdY9ByVzHjENqSYyx
rsdcm40LYQGTRhNa7OW6R9NhQ9qdgN6uXwsrFEV9/TJUZ/fgPRppWoAytBiRJxu9hzNbdC7/2nVt
RqfBUbPtBzCZbqxPQunQlxmal09aCxiy3u5AMcNCRLLEbyGgn6mLH+93xKM6wn4KFSBEVE1KZzqE
4qVcee2Yj/sERwnkASQ4ZxXYRxX22ouAyEZYaC02X5cDNcec3yaCH0TuF257W7moD9TIZVd8SNXF
+agQf0Rn9NoTvNOsUe2SgLj2+ZWnzb0BObO9wOjbcOevSLIobUV42elADw5CR+0GNiaM7ECTcAbO
kMpREDb991XHjEPoNom3rBLF0ymvG51xCUXhg+x9a8C+rkydDwLvkAEo3eO3zijPK7MO7MyWXvoF
eRbVKBKkQIOvQHOsj7hbne7HYSzl2S5HzOyS37NskSEWPVbqLxAo5QhnjFKKliRiQAe1NIX7mzTr
l9CDWqcMrPnmQR/AZT3YYRpgtrWslL8iPN6F97cvMyRQwAYKL0lPb33/BdYnLs8yQjrHu0saKTZA
NcbvIJQSF/Bo4Tu8MIsZZmmX1I7OTK3FSl/rLaSk3NIsm7KCMUVmdnwUF+yqSx90WtU+ANQzQJqv
m9yk/gTHUZN/mhXusN3DNhmP3x41ZshHY+DzBS34y0RCwc3P3mHa4SIpnEHyJwmswDYTbHhWiYwv
546YZgDfenUZ3Vza/b0mKfkmaWX21AA91TQBhOHNLjGZ+4riVuD+5xUFYJ54beCwRrswXB8vbUDH
lVlwVBFfHIodQeNUjNMqHOm0xd6ueompqK45vqwUxHKotFMk2XJteqZp+GA3h1+g0YPGPKC+4fRU
j6HdKJWBJGJjXBpTH2hhjsq8/g5iqmTBpMNuj0MLdbnGdHne0RTmXWpqdBEgAiv24pyR5DCX8Tdh
xAck7AWI726YUySoNMg2y+HKXp/HUKJt7umzgB3OHrxw5dtOrLCIgD6eaBJ6p60KGUUa/FruQybB
OwZIY6w/AjEyBAOm3FUmBs+viA0KD/OtK+8erMVePTYoSvII8kQ30RufdabbYK0xS2/KCbB41NF4
FD2cX19tWpEkUeswCg27PQPEJNmmNNXIpcuVHK+Il6YYvyWA35gdcUZZqQs/kwGHjwwFwIXuOBeI
WhgkHREqBRRlcZ/VT6t9qBidQo3VIiObpEQq1fIUijHgWs6TXAIxgGopmrzoyiU+GBxhEn9VQxv3
gwGxE2roY2nB4z5RoajqPLk/V30pnJSIGpChDY+D8m4uUbY2T+pZqFuv0L3MTbbXYjgDqPuJR9Yf
Ss0psOTl4VMNVtxReduFuikGdrAzrsEMcbXG30zEh0UQnjZt9ZMPuDOt58S9iFHXhQkc7xGlru18
1DF98tXfnZ2xCPhJzeiVGpo5MvJ4AyWcKdw/D8uTG3vIYHo94F83a48Z8rJisjXjBfkVzdogUDUk
LZ7e4GgahiFuJMO1pxKJDNPJVmIQ77Gc8Cbjp16MoL8t/gaSCumsriBpIxl0VQtYK71yAbR9Kz1n
RuK65K1YC/icIZfYF3yvYGvWWmssmWwouMPbzTukiw7A4O39iWyfE8ME2UU76w5pCh4KdGj6KZ6t
deYZhYhK/anUMYBBUZhSbfnor3noQMiZSHAvVqunc4N5UqlPfbGhh6mOcAeWb/0snip8anBhxcjh
GVNJtjTfi9c6gs9smHPJemPGq6JDnvGlhdB+gplw7KiQLjmgRwzSK25rEmZWLf9nhYsU7/+ft341
JvEvt2tzDrBLhgyHBjvK8rTBU6is4PCU8nVi6795FXYkj557zhuqR3TSID0nuo/PXB0e87jgTeVy
0iUiDbMjKC2rhPvKbBgzdk9fEKIVzBVUGEFv9NRCywZ+y8Cv32u04RnA6e2oyMlioZX64ffUcKBy
7NHUr3oz4QD5WBQa16jXVeQ349cbDvLLn/UAc5I+Lr9aokC1anodNqXG2pIMKW1oGdjlS29oIkjN
Rbv2/4hsyEWWz1n8vdWK+1/7vqEGV5KidgNoKwxiCYd/D+xMEoH/Jm2JWumg8d44OOOWoJaWCTbp
oQQ8OiF6v4wZAhfmRrxYNoX0n35Uh7qdwFB4F+/duuUnT1p51crLvYQH/aPS75TJEUzGWp1pnt2w
ew2eGYMnRBPzMNUQGtBfvVn1IZqWZdpYs02MxfYtT1QPCnF0uNaiZyCXbMMr0dN8gezm47ywo1hU
wbFSO576r+ouPTqzgGY033gXsM9bM7drPO3Br6nG1DlZlXGeGpeOVYUXBwY9BIAA7TXMAG/qj6mn
pop8M2063pb5lPR2ndEFmyynJfD3C5adNSoY/AARmiAr35cOG5Nv9pVtAu6fe366MJogLj5Z/fPw
WYhKF1Rhhj7CsTxHvhdLp/PsFNVC621IITsot3lgfwuzERKRxz6EIJymlcE0JwApxNpqxaVhz8dA
aKU4jQXsH1504wEtaWT90wnFpoBkXEb5LcPZcoH5mMrfT82FZUL4ZVxlnNbbosqr9gtxJ+jfkYq5
xUNWjAx9WiUKGMuR1ReYkxTXsTJC2Sr953miqEHgpoGr3JBBd5h9MXfUr3yS0zfQ9qdyeU680dRD
5hyELOHGrAk4FiKlBQ8l2LNd/BqdjQF3DdwLezDmfLlfmmBdvmfTqxGQMWfBzezgQqxT5nG9me4d
MmtzobuYlSS3XeQYC394te0sX26C9xfG/ritR0nL0/NZN4IdaaATR4gQTga7r4MLRzOdPXwgPyzk
SWvrIpdyZwhjRLH+rQ3khk7U3pwfMjvrc7JHzkwD+IeKFPVXGCTod/9lXlfxAsVz+GdJResJWdiW
SdZ49EuTXduZBUzxQGUt3wpdvNQ+8l5fl4pS4u2aByGjyXWLv+JNK+EVJGy+SNMNtPvbrvrs6ahG
vlHyDP5COLLN44WDm17lNqjnyBRulVkgu99xo1HFIr/pmO2uCQKVygHsn/YduIVDJXlFGpozNxI6
SV2HSUzXuNohPpv35WOIcWClndqeEhAGolE7sG3TcwXJ5d5ilJ3IZn3bqobypIEHMWoNv7BzwJIF
PBsQCFBGtctURWL4GzUaar4zuW9rXtHx772jOYE6B5+NR/9XpNrgfzk5xdo6xQyihbWZ4qw9oVK9
J96Vb2suwAn33vxql7eY92cQVTWcMupm4U9qgMOKns9HCN+M35ZlBnA6nHP6cfuEPcnnyToPk8+/
pKxP76R4K7xaZmYG3vWA/B1NkDbqw1e1M2AVP0SYt5wEHmfIxtyvTfq6VMlq5EJoLJ921HLo4abK
lXZe2EoNz004TW3BNjcQ7vihSF+w1l391s+86QlpluG/ZI4LXdIbJ/V7AafLOO9hqY05mShkWJVm
1k53R+nu8bhqKrnK74tEno38MsQVoNHWY6Q5bnQB+ECqoXrsl4+YgcznC+dWT1a2YawI/fvhYKYA
njEX4YihEx06uC0nmcKeRhTkDVa9OrVipQ/LS+4RRqGYtW42mUiLDdz6nzAXYyyUF2lkFBKunitm
8QqwW6EI8XdXz1ZoKjPTYfXrF+S0fEpLLtNTnCHohe/nHZVZ7YKG26lNLIEk1R83MiM/vBmBb8hf
wBaFShAem/KyAImokgMA7pSHvknrFMfwG5pk31t+bYQNanhmlnl2dm2bsZ9v3gFU7UgUQlbRWLAn
qEEGKltcD8WNJJ94tQxCMHk6+jPcXmt9cdNS/o5ainnBX/p6/Q2KV0lNN7zyYEy3w/TPeUqY8yq9
y4D0P/uEddf/22MAAqXL59SLNhPeA+ifILd78cC4fxbcai/zq8VHo5fSP1ottoYJ59MQtFlYoyGi
yB3Cf9xfrAZS3PlVTYlkrBdxCb+1GFGGesdvVNI8ZcygnI5gJ4REz0+dhHcUZBzPWsl38H5oPqD/
KTAg6bVgnYHpF4BVJBdE6p2VLNc5oViRh3EO1p6jACK8FKuijTbNDO6HxSSzDnDb6RdXX/JHy41V
icNqvbZKx2pW/+pKsoCoElWwgVEFgKkjZA3hFakqvDv8Y0ONIoaIdClyBdaNPQE7mkceRGPQyY0I
hobJNW9jnBkoBeYFXwdTFOFxhicF62oyXlZCDWstE5KY62irQzglr7DbeqybGeHnnzBfkuY9azac
a7yVKvZpNzRl7ECIiiqYaRKX1Dgq59/7ybFhYl65HX/gjcJpOFo5V1iTslMMLwU5Z7GLV4uqMOOr
ZdS5hL/mbE/SkZfNOK27bc98RdT5thoYjEzz7CKfO5qQ5ntFWEbDIaSXUO4lcaVeK3b59aBTgh1Z
UUGLjoZ91lqV3VdegVjv9b0hdwchcLR2t3C9zL1qJ61zMRucmlb5x2WZHvmI7qfGx6ixZsHRdERR
L78wmeqBxEwAvzNHwwwGZqooHMMcGXSJXyShy4QW3IWcFkK3lrtR9Fsl2Qbl1Go/vLfnZ+n8bmel
azFGBMjZFMZebZze3GCKO2HrfZ7jigYjspmQ9f65SFZnEMtY/EnzsGA+yPg8mdNpKU/PTaCqB4Ul
p5VwO+tqUUaiC7as17Qb4DnNtDE00aOviY2X2QprOdv9UcFOnDpKuvUKCS0YbT9LMtlHstYjHs7w
CpIBH9FpmLSPedlN1h+8VNwzpVvNT3S+Vqy8JoATa2P0qvTYv0lrBnBy52IsiLCUZf4IGKHyUup+
VlsYdHhPecK9pQhXXjqGsrhyeAXKO1Z5r1bKcOWmrCOzzXhyifNoKbVBQbF0aF2cPwMhr4IHnfTL
BBtlM6e55pNx8qhlzKpkK/7yH8PnWHYV52sjhJMGfHak1FL0DzvQ6Z7P76VhfzeRM0FfhB/yRNW/
1sv+QscTTq3uG869Hom/QEjmZtEbpAr/SpUZKDc6YSO0fqL/Rk8zxGJvCc/HK/swedi/htgqmJe8
RUINj0Aj0VCRAe9NCq1WI5fJ4Ca/R6vI/ghIZqyMd2ncPGMn4QmMMVqQDBVD82fQ95UhxrhqxA6A
W8MIhalvoRcl2Yy17JyEWJXlkz08pzn3VrXF7dvPGZ3Kl/zBBj1SW/O7aubcDgBvpQp6PkORVVpG
GFwTRmyGC2RTSBRmUoH1bmZCsaD2QYJo2Iz9iLhhzL/J+p+inRKcNO3QJO1UfDmw4pyUunbFLAVT
zGCC+9i5a+5l4meGLQGRdwFWpw/cuB4gLDfcADUkSAT0HSaj7QrE7eEOR0QG7NSNJfuXZE4kO6NC
nn1eqQBlJ/TtOgrR/Bft5vaJ+7MPkfOPmbpn2bEhSRGeNf38h8qH8I+NeTldqQeUKFw6dX0oP0Ky
13nyvwoyEqhWvMaS2fMsjDrY6W4Dr/0jRT5d0cEZMUxPSWH37HK4A/ErO5mE5hQAXxrMKFFs4kn+
3u9oqlNU1l1xqQ+aeOb6SU/NsxUDBI0cRh3mTfHFixAnNfrJoPqTA0JPLgH3SXTWKUauQro/z0Uu
cDyMipxOAGm3D0AosMaqDIFsYhVFxoaKLSx7H/356vNtlErRRpmMWjmM/MaWu7JHtdmlZsnuAydm
g4ZK2btdAYwqdVYa3LikvNgQobDSeorRB9tnHzgyYRRbv4mMeCsEOpTxEC8nAQB8NzQPi5XzGvI3
2Xsye7WXpTGZp1TWbWtbPLVieS7xZ61iYLrRUtM8enXX0oywaWNrp70TbsRqSFSDr9kMUgrLLppp
GMj4mWdGNLhAXMcoWfCpAfUTqghkWO8KTApyD06VOzlBoHprqqj1P7gp2wy/5ZqCwGd2WG3m7z6E
fNLivGy2c1XxhftzLOFPw6B/CQijKOiqUZ7jzL+q2hbyQRm7XPf9shpuNEBZeyTX8O3pAO6f8PJ+
CW6AUQtrKWRjWaXBvsE7IsvMLbVQM+h4KiyPf1MBro2IJP94KwL5nxNqcF1V56sQ36UZefVl/hMR
+i4rimnwANvDy2mFFxYD77TGO3axfvRX83Z7y/Jlm9026NxBI5ls9LusCFrEGyCBFjsIYs+1vG3I
MV7jLNkqk9Eobf90KCbNt6tzZPYxVPXZ+N/ROYjZi3EQBpNHoMrRkCntCEgVajqZqhtA3rok5ddk
g870GEMzU7acBbGQV3Z5UARFgb5jxle/qubDHDyW2Vu68e9Fi+DFynaeX9IjJxQBqMkeHirAENZV
SabEeR7fFeVYpy351dg7wuvyc+6GHq9rB8AZcewspsmjzGaZXTGYZuEgyk8y8Pxcn4WPi49PsA5s
n9D2jqFV1FKK0Wrx4lgiomtXWqJ+g8xfVupo8xCkcb4wKjXjS6gUjEiGsM9i21nHBnnEiFt3J8jD
CZQIL31c1mjEp3hMBI0mGUegUIh7oUJx/uCFojDvw4x7PgDTt+28RUYamWEnOI+8+9reROWVvcqv
YqsVa0FQsT0WX389TeXMm9gslasChUVv4hHM2mUR0rPhJxHWmKlApqG4aUhqsRfrxziiqX7x6Tgy
7KEJTb7eNnslTLP24aIjfPAgkMGTJ7DgjYMRwm4OG3LezfMi8fuBX3rMj8d/ynEJe8toLE7RbPUm
lI4ILvvr3m/oHeprCQd6W4cXvWRmJdgF2vBSmiMHE8pfTOOqrv2Utx/myCIWdI3ONW0LK/yFrSk0
MBfu9rv63XgdTi3KFaGXPZPhA8IRd0CP9gqDkJC5Eaxn4poMBrA2H8xgxb2E8UHjp1cvKsf4hm8Z
snNRIpDo6yFn/u8sZFRvDzWS8NYzDFvaj4odr/DqP8rxDSLKXsDs7XoeIhkK81L16zjC4sVkoW5z
J56XhaB6HvfusOzBL2k9vQX3YAKcLjTqyxE0XOrrgHDr1wU1noW+62Ejo1dNUoNfP+OQExQu/S9N
jITvKRnsmOwnKkcdEQUWuOjitVOkRASUJZeNi2m1J7ILJL+XJpxwAs2ZB0KtGjQQUeCaX0IzCmsP
qbLD+64v2wZLk9N85CzqnhA/PyciNFCHKDxqkv3FBI9dXo8W3TK14Ikt+3VAVHuO0mVoBTBIi75m
rxUkH0Q9PEOgKD3/rgswsTbOd0094gC3euov00cFMye+bENA7ahougVvA1SpBLUzq8FU/93q1RPP
0h7hq0PMzwvuuKmF1d7/UF2jkKvlWTTfUJhs6ovsNYjD4hzw1hf9t8lPqQTGryKmUXluRXY3XD02
f7NPckqG8/qHfh8N4tNgftuq7oXXU0quAi6WsIBERZBlLPU9J7RdC55yfhbvzxZFHE9R+OIpBpcT
AolPtMGViBC26ofLN38Y3hq/4ezFkMqMbH3YXMrFb9FoCobbbFb067R/QAh8wrfnvlwXeXcGpsr0
9rtwaX9ypr8hQQeVFB/G8qTDMNPi166HZRToS52zaHTexbOBRyo8+STN1h5GZp5/sFE8zdbYWwge
RZfDYqaAMZCgvSzu+1XdIeOuu8gDsrWfn9T93TAazxxyRAZfMwAoOVtSfoL/EEDG8sHe9ftKM4yZ
8qQL0hZ39oG74uljvX+CIY62XzfGrOfXlo36ESsHZAcqGEuLtWSGlHAbbmXmAHMO4kqWdEulwLq2
5f05cXurlKNxvR3ONCUoJpzGHlvYQpa2h/zjxA27q/DS2rHXxHQNANC4yaAk0RYCmzLPArHFRpLC
nAZakYLUAAOZyKCkt/YVpPcXxQpf20hu+g3iZu0+vj3u3VYTaZnZqCqq3iiqLxrUaNTfqN2oD0rh
kmupNbeqNSUd0xOWlDCz5R7u0KqgCinWH16oeetWS/mCNV1XqGRmp4a6IRgpbEQzxrDjLnEaBs13
ypHAU+afcgtockt7Zcw/462WCkZEnjAYkASAdfIXldH7HjklPfA3r65fUFU5ZAzQNKji0NkIWxvK
qhcu907YUo6xz8ibLKxSUpe+Lqkr5iZVdrMjCO+WX9poRdMDeIJrWm4bwLLMxf+bEJOhk2pVG0Cd
4UhokgOZadOHKEwRBZpO1fP9UEC6zY41ImByilM+nfjncFJStn8VfCEvwzpwDqofKk+Xs9whrvby
fgeNdTkIV9opuznCJviFl+MMIwKDNdQEWH9gql138gez7ZMq7y+iDOwCIfB//0iH6xzojwrC1rjy
t6Ip58rCG+B43+8KAIQ1wh2ZFZsVxOFZ7uKXqYINkl9sgOPcbF7nWsUOCaYErveGg5ANk84dDLvr
UitMAcoZ5L24Nz1dliruYSgSrwFzBz4tvdBToOF41iW0gqMEKmSADQ/lItUFNUlm/OkyuRl0KieX
VuV1z4mGFJZXuFjHjhLukoDcxxjTndPLdF1hzscSRwiDbkq3IZ7AyDTYB+fyMIPI4qZxkB42E7qd
/oFKv5HRfRatE8TPVvdmTcD5jxTSxiAFpyVabxOj/J+VHEYG59FM4s6tPfmXf9dvyKn9X9tG8DK3
pi8OwyUDntuxPgRorS5O8wpoofNXpR/2rBQ9U5JMSpbA6YWhTpvJPt71NXCseH9x4/AxxxHAVekP
ojClBE0BFgZxRiaRrEL1omd+yNkRxGYVI5z65Kjqr9aKbiQk9HLGalroAItT8mr0TboUinsq0Z+3
9YgyYEjBc1Kj0qw19ML1Wk9cDszDXtLLPOV3sa17wdQLsI0mNd+1E7ZJak1Vd8dIRIuEzVWuVny2
86Lfe0K+jgaatFCdp26+T3NsaCjfyGysQ41KMDlLRVhocC1o2Xw4qRxTfYehr3O7dJ9mowujXniJ
ZsgwLqC/7QpCbU3VN6mBNb9tEJ3mCDsLaeajQxNK3LeB4KhYVrPfACqjo+BIWrpsmbkkwFdjV/cI
T9uu7Q3Wf803pkh1Of+qMDTGUklqe7DgDjocwxuyN4SkBce8ImZKUmyrPQIE/75DqRx5SEbP/ZiP
OnTI/R6RdGzyRZsXIxgmbCN2Gn/GhJ3pweVEoBzCEAga1HPCuB+Wq20eyC55dP4JpQ3qh9lbG0qX
qW2eMwUT9pyRMRdoP5j+E0JFdS8eW7vMY2fh3BxjloP78UjIxaFI0AlIDmYEZowM/F5VTn9NRG/q
+yIxBDzrUCX/88fx+WtLFllNcetPW/J3MreCg0vkl9MmwwtcV6aHIjaelW1kVWwJ8gNjcNb9gCbW
2HllehZHp7NphyvhUBfoA82bSnGz6NzaxozAYzBzcFyVN89lUrzbPr+Jb68ey6PxxZH7/I5W6tnX
3SV4qpk4tkWPrXKC9Z42ecp1DWZ0DW8VbieYOVwPZ8aTB9YQp+wCLSZTgIONc5ja70KQaFuknznU
YGJFG9w0+NdiuvemGcV8l2elOnpmYBDbUW1pN0nKYOBVECRq+Cia5sTSql4kb68hKCf0S/FUe1BT
oGusY9AwnZT/yS5t/kfawie+eN4OTXHb41H2kufGpNGg6lGJxWeh36qeZODg0PmAPduWeoKmeFtZ
zGePzjNZBFDrmgsmaBHGQhhtKm8Po4GIkhQ992+UQY30h/Mq/vIwUkwkX5YXdM1T4E3eIbTZESnv
Lxa9QkV1jGzlIu7UyqOAIGb7ruEW7Rty0zYs5tavDouWjxVOHBEmbW4uH67PfxYamMkF6rwYklrh
byEUtJOhuBboTUV3h8R+zx9b/zQo1navzXxM1vflZ1rqAQUpBzl/RHqXQfCjc6u4UzIN+R31F2R3
z9ORYJGYUmy/TVeAu5t6mWu/hhs13D9IdxoFE+H7jVZ7ewcTFGlMdu3ZkWsC5gr4RQyrXXjAmZe5
WYBtpy6tHQrN+kkC7EVHhaIaRD3gqABwwi8ugHExK8DcCdruYAuXsIhxu4Uex/4skidY2ZbqTByR
VRY8hBCC+H9T+Lc0zr/nTVdNwVKNpMfu6fh4lkzpkT+gdk73ykxX77Ksn/IhXvb2ujoTzynTOrHX
Q4npDmkeYDZUy4sgZqsTyoyhOoBvmONt4l7Q8uucCtAEtvugt2YDQK7vaUrhPjgv+DXoA4ifRhmw
n4c7jtoz2q1Nuup5Vi145BiG4X/+ljHJaFNe4tUeTVHxpx/jxMiCXQCERjTBA9ObN9mmx+jBY5wP
PoCA3kFKg9vLon0YXibECZOK8e1Lv/gJJGm0itlK5gZPsMlxhckdxyKxveeSjlQYCvcIhVblQAPC
lnJS3EXm7KfWRwW686Pp85KcAok/ifuthIN5tw2B5d5yUSdlooZk8EohjeYE3z5lc9yUGSiToVyl
Y8ZkLcFe1HGPlhuZA6UyThBbQi/az18qP3Rt3fyrjbyYqgdY3fLilQJbu4yaV1Iy6PKe8rRo4YFk
f4GckD0DhfJCvN++j+JcaolEsFhZXwRl9ZQAXwvzYGq4OCMarjY1RbfKvFM7/OT0JYO2uPa2LPd6
Ndq1dn91eoITC0A7CoaHt4flPct+RcxXAKg8oaOzizUOZG1prkscGi50nSCXuWLYT3hTPnWxwluE
8HcxuAYG8RUatu3G6C/LUTpHA5d94d9qXlShUpewJCpGcHRqjEihyPovTTaePSSs89N2J2YlXHjr
DogPAnyDr4tF+EDav51JF7Wq94X1amOKKDntUEeSbOZWndDefjnlgADxQ7Q3WNSXfQJSTbtDbF6v
SWDVWOIYSrWtuNgYXeAh+dKEdI3DTy6Zwwzy9jmeG6PkRvbdXwbp+eR478k40SeVEudi4Ur0W6wI
7aRTvXGT2ZqYpKprLuF8jfyrB+UQWM2PPt9GgI6/4WiaNGmWmCf8H8twfZf4pLm1IqWyEVDaDkgf
mBNsP0pRlbT1qnV3+8bTzc1QMfhu8ZjziYncJDeNWivLzxGiSO6piyCOf3KaNAi/ssGUfZYHvAMT
breUM+xYtXdvECD1OxowGXVfVjNcj0lxUbxXgZhjuHGnUu8Gzrt2ColM4ETMWwxezivaK7F2xdvP
YKbtwVlEeE4NCDlKQ6cLD9l2M+RUa75c5ZcuElubExVu0ahRoXqwO/m/lQ7IsA4o3Nm96f9o4d+4
4OhNy27YSrHwT8XNjvy8AZzzMmfBxt/w+0l31JkJIXYubhQ+b+5NBV6DkFv2F7jN8fdMR472+Jjq
yta92v/YJ0mgzoam2eBxDBMEXzY12oGc8BsOxs/5HrbYVA8OIOFYIhN0aXIhKjHz4xBxpRWrHda+
QkjEAFTeLF2oKobOmhSGjR8UnYWFwZ3IC1AGZ9GBlw83NQcGupqEb36zajxqQMBV30EV1iAJENu2
So1WxmAgLqFxXscYluwRnw840JxPJ6bHJru2FciD2zCiUeav2O5yMowv6pnPbtgfJuzgngQ4+6nY
QatOt4YbVW4PNkI9TvBtHHHQaNcoVR17pZv1Dp3YMsFhxfpCJ501AbR1sTjHLFegMkZIgAhc8G/D
nZ9NxhmoIFnDh+j+9Pnm7BYPI4Vck/dRhJ+0XTIN1w8amEB0Y9ubEzvozJ2Bdirb4EYtF6pmLuKg
UW5BgZ9V+GfCsvXNDPYdwSpRabxxXTqLj3AzaiQtVm+9OfC+DH3oKCahZVftUQYEcx1CN/Ah3FMq
dYMU+fRsp5X9EqPsCB3XYUimmqen6MQjyz1UrDZhHwc0WGoXZcXG6IlaRrThU9uMsdAIYBz4gFMA
dt1co2E245bZI+xtL9u4Oo95fGDNm5SMaopE2CyGwinmQhs5OprwkWejNNG/9S0u0nHFJlEL93td
2FEm0JAXz3aAPyZN6HD9TPC6h7GDepOpFlnDx0VHzFnhvMFKOtN53yumPbCXn/MezAuBwGfAas94
rhOfZ/mqV7krRY92RpfqZFz2k3/bpgKnOFEJIMbzQsmld+PyoIgDRnIbbWOZXiREV575Ckx7OJrF
1D8zfeU3QLVxpbdY2v8nGj6jyjaE7BoMqopSaM8K/Qw9eEltVa/lbsy7OYgAJCVpt63IdnrMa1cr
RMYh8gPNQBhIElhCwmD6a+W/BDm2ySkPBq0F6amQksI8hELz1zU66GUVF9A/n03YZhaH40XqPQOM
fWYc2gLSXdUJctPa7eTEH2PhRurNEvGTil6EM+dZHK+X9QflU4k0/Fe+D+BnPddNL5z938/k/2nC
nMCmZGD9Ws82adV8bKa+B/ZhehJj5uId801yMWNx4i2wp+ZGVyfc1ZT8j9mIlbhaZmyzIblAM4MD
l9MOfIvXVbf5DLs8EJg1qPdNS4EQa9iO1GlrUJyT+APWdd+OY/7zwbutbog6qtlCxFW9AftFQ3ai
1w8ZDyoPFeAM0W+GdSFraNbdnw9OyrSd203qFoJVduepBuW8jQ8px1YsBVrIy3PpdUUjutgFBBbS
IF1zBx6F/EWo2MbKOr/H1KgKRL4opeooRei0RfdIadqc50iAhe8eWWu9bkEqTsMnWuMEAEMe9G6O
RHnxzsKuk5DfmzPfNvGqxAGlbjdbGyZVCaUf51AOxcZPIf3a2F7JG5K+VRRdXWWs+2xq8SnKKxvz
F1KjPVYaXLN6ZKfMzPBvaHZCFrxVg1IuaXQeYWO0QP3JfJV22FMn6COBJ++Te1kPsxXFVlcm1k8x
58JJ/U4b6S2h+0XETezSzHreohWSuIMSN2HsHZwCCYaLksX5/3uQEAWvPlX3XhgZoyEFcDchUAtu
2sC/41s29EXq4cbuIgbI6M5lSxpGIWGLBZlQNDF0KBJDV2gHTr7Xy3HNUKYwvF8+OgyCRYYdCF15
AsVj7XBes8PbyveL3s1cnADF35hzBXrfOGxWupnIgoqWSehG2SUVPeTWEinN/daMKTnmjMRnxGpn
z9y2MjjlrWNVpF6aO5YHG6WWuXdgSDIH3JWcRNX7Gh2fDhPS8HOMSXLagPIXADEn0jNbGU9aWo82
t+iw7jatkejRkq1FquEQ2fyNpm5EgLKwOTP2lDePVpUrZ9IPQetEm+3QktjmaS8LdIHvEoHnuPwl
7kHX9uKG8SHLTrFt0E3JjRUtYJanT5eXOhHGoi3XFL5y+w5Bp8/SN0rnFizGVUBWstpxlnOlDIrP
tOk14RZP7/HdfcahrLOJrxGa8Xd0Y7sNtB/jhTvoujy2L+NgcPtTSouquHI8Z6jociRbPmQKaMgX
w8Z1nxUys6S3vMYlgf6ePmc3H6kSTv0HNbT7aYV1KzCfkYEQXMyX0EnOxbC/awd3SHXdgYo/Ju24
cbAGWPULArFoEq/i4zN58yRrzQ69nYXmWR06p0PfCxRUiudoSkvz7pbiuJKMlUlMFMDykwAvID4c
3uAIGUDWx8+uyTRegxAfoR+fyiNZy/+0JOGOLAiVOWTkqm9Pci7IEMhGjvOgxPahaqJ73kAPjsJh
qQT3x/K21RI9S5MsRqmRy/Fn6OrHpxM/2yFusJFi+ogqco/z+Ei2gxJ7AgU9Heu76KcM/iAkZH+i
sOId5J+sCUmalIdcwAWy47FzYKh+Gdw8havpwCKyaOakpkgq4EhDloNpK1KV5zuJQzb1nNKtIass
yWxGK3CUAsWpo5YTZhMmH6iU2xDtCXOWqcoRjF2aZbvEPmy/anDLScYWp5fw9B6ylXQSQ678wYVt
UaKcZT50Fdth3eGmQoVy8lxjf8ApwehUsPGOZuEJLo6PFaYhRWXaRjU6ozQVQHcrcagoKMQ/9HL0
2m3IX/GY63Wnu85lonY2FjLCUT7f8aX5DjwdkmZ1aKMLYLWuf4IQQahs17WokvfL99ZvHN32aM8k
MAlONSb+m305otbf8HXIJTUwfcuVlpEwkBfewWDkxvNxLl75L9BcT5f0XtLQ1R+HSaSqKWHZv8OI
wUihYu9AzqgO+e9VzcVXcLJDgDtm7DPob3Q98vNMsg37rL54iiQUhACmc/wvnnQvuvGyLBdL63X4
aijN45X3coukDgx5Gyl35kh9jru8AD4lLU7HC6aoVBdaT4GzsoB4uKhTBoyGQabRKwznHZzBFNBM
lDv53DJizR636T59cCehZd3/0Yydaf1fITSZwWwOYN4JT4V0+3I9XMHINE/CCCJB8wLJ1XP8HEZ1
OXTBcvawQ9t8bxN2oqq+8ux6rgZPUHhkPfVr+55VpkTBLu4k3tg02OF9OoQRcTYlpEqCRm1uyouO
WBvMRoyNeZJEB2CW9140FV9ibDt2jKFL/UhLZKN678fOBfFmtVdxGfJ1tGli+KAjfToPUpo6sCyS
JM/GrN0UktjpfzHt9PytHnqytnQomDln63lN4uBPXydOMEbD2vsFAv+rtzRgLrFyqnc9IM6Uqy0r
Axs3rh8c7x+4eL7O4Z4e+y4jEbse8oz04w0U+XE+ytQaectnR4SKf3dfN5lJvjAsky29AVFCUA20
R1hZqS8+6utoHOZMz/2xQBl2/RQcLdn/unmbwRl0RKQxdnkd3arxyNUUnRuDcN7AqdzeciAgqEy4
HLIJEPDHq2n/LUylXuSmylgumhevAqwOKT5JlzzfJ3hkmXZpD8c3SCxtaLws/e4u91S/nASyYydh
GpyjgJMsFgDfgTc9RMr0RyBjA8AotxLjqp+iHsxqvwlLUoA8itTv5JmzonXoaePnHlUykIrJwGYc
ZrBCjMlrnNrOzf5Jmb/UTDtphY3ji0DmdyMm4u9QgTjAdUY0ZiFDIvgTI6v64wxbqTzZKask+ZGs
771LSjBt+bIPxwscfT+tMfoA8biQ5KxG0Z+iToYmWHzPFn1iy1YPEY3qMvtGNKD3fD6lNFavR5AL
XiV4CAqZe5fURXezRozkTMFzqkjuamxdyuWF7K1HOgAL52VTkw23n//RbPpS4R+CcA8LR1ziZlaR
o/oc0QUBiT/Dwd2ePJyikJJydN+IgbbSJIN51bOBAIo4XHzgIH74JIgn2SjVYJ87/GQv6P1Klsou
JPPtnqQ2a3u4tXOhN82heMUps22627dEwxSTfEpUKGyerWpmpJSY2LiCLWv7/kaOE2z1yyvkgt56
MBTtIcJwrTAKaAzhB1zEQTeyGjqb52WbhUAgPId8mRQMAn7syZ2kyCnCzvuH2YxB9oRicwmK7Rf+
CujLoNVPjgd5HK6wTa14GJZP7MwR0Ol1Ojl2QWMS8tjX/5YiJde/y6TUrI78JEJ3O3qbc+LnfnW7
9oMk1KU9YzunFSQ8KCYv92GHIwq0By4zQ+D43snCGmn+7SYepL7GNV9aI9B9rodHewHVhOUFrsjB
S0etfMcmhaAgvpO5KnK4ZcHMMAu33Oh1xeVH4OCp0NcsbLxh1/DR9+ffWH32Ju766q7anrwqerPh
xJYM7DOHddtLkLNo3f9MVsC1b3s4k1IKociKGkBH4NAij6Y3+f9wgoq+cMK5rwGPBa+BPvkLC5d6
Hyn32YbRj7dMY5xlAfhb+hy5QyGt7USsmKiJxJldKHaOODbv6O6jX6/Ur6+Xzvoe6qHSCf2RmJZU
ccdoW4Ngx0JpoeJDP6G0TQ0+FE3q0bU6fB5KaBAvTleTFs3bS1qirQlLHToC/WOmRQX8g9wrvsnq
3EBgJLMRnNqQVUQUBOovCWq35/8ivsuW8W0f50fC90dtkQ3Vodfb5yiVM11GBqOk3gsBGrJ7z2Ej
xHQ386TYrONnbyxhSyPiFOkTVJNgYQCCiErWneJkOR11t0X10yCX82gvrtNcPOO05ykhyLZZJqUI
1JVYQIZxzhfAWhgKP/+IR/9LR6HMPrsYYBAV3iTJg85Ilp2ZF3ssro/pHWtP+YjvctufSr0sNlRR
oz7KH/3eWUYrEkMmHeVbWfK6Zda5CeLlKy2+LUpkebnRGHjsWpv7tMhKtxx0DT6otXMAuZni7E+h
9F9qLCXDUll60ZScdyWI3ae51VNidlxxpG25d0DZ7ozEafE75YaEP3xvuPmkkjjopbQbkqW6Um+r
FGkIwck2MMmV6j7vsFsz2Hsgy9eiwwUQaVuuT56V2sAWZZyEZD6oKl3qtOTyvwClF7EzLe0ox9VX
5kdiY0uY/AF/5fskNZqNo4BfoObJViwOEH2HjhJ6oUeFiWLSbRervSPZ01dbwlJXOIPVgX1B8879
sDn7JugZ4Ca4vfXFyTFrEcwcJcZuVKbZbojQlfLS2RQKolyfbbEVKW7eagU+En3tXEfeXqmfbqKp
/GgG4C4HQYrGzRCsPIWO+8so2IgNbyNw80xPTIQ/92vXJ22syEw59Zbhug8Rr95OD9Ie/HkjuDbg
WlSmyrv3xFWavXMWRzBSz1ypybEa3Xt5ZIfdUeW7JxbgbpEV+UnGjx/iyydjgU8aN/RFZdMjPGU4
VRFXncUvTqkZowvGBDcnP6cfBOWAFV8T/xlMc2drg1vMu1DcV5wzgilp3tbQKSTk1vOWrd0OO6ps
7SWUCV4tQiEd9Oz+AwX1uOZP4UoCOyiWOr81gCM/Al28fD3KK6Y8/LpvnaVK3Y5aieKyzB7hgFZn
LyMYlIJ7ZYrF5LBOOkcLjw1zBGdYHnrn4xB2drdngMwagj0vNVEllviTT5rWsAuQ/OeREK0R5lsQ
s8WiiMOjPpEdLzs8IbUxPJSMlZf7T+M6AuquYECVYEiV/eDCJskeLrYrylpvxJ9vF+rA03VRtQiV
2QxwR6HNyxSV+3oIQlBzEAidKj1+0VcWq9Qpe7veqjZ+gfb9MkxykZ5Y8sbw5iYz8nvsjhlHld4v
WiG/9+GbV7Glr0Bk74g7a57P/YMV/nYZE01V47KsyFkXniHCtK1OnybC/I9q6lvawAE4cJSWfS8C
wrQYtwdkuDMy7p8ixhxBt7kfRvqsf4pbX09jSGU2BOAj8T+TY5bvLwKvrrYdpxDH/bKefotxnrRc
rAS9bD+cp7vL8QpCJCj+A2lRCpNfAtj7KNOFMUnuIt2Hi7S9nsviemsNVkIcjioEPKKR1qQV2Eij
O4B5627ciiHfXkyaVSClwbaZzmVlML9j7DOSwUeL6ZRXysgqE6AYH7p1hWI63JQ6dJr09zuy89kW
0i2xlY5pE8Th7q9EzfoVbie2eFmfdmByA06cHMuKKBwxr5dSIur1KMEmrImHiSGWa7jsbQlpsQVr
A0q4ADXd3TMDamUvojoU+VlfkgY3OJ1Ny1e1Z6njrhLPhL9MVf6hmK+4KPkwSUnAmD3GFmZe/dAr
LbPrm+H/aPmKgYu91z0Ua2/nTTQYMjqhStyAz5yikbAS9NGryaU6WaNPVbUk1sZU4yR4xxnHkxJF
DtneTQPUi5VGspd1G1PMevN27YkAHJXBRgFJSe94PBR/QJ6cVhu3EPWsi9QPSRLl1rgSS5kVJLTd
Bnf1xO3/Sv0xw0DFap5jt/VofUKzVV1kvVbll881/sGGg5F6emukFiOXTtVKM3zr63y0zG5DaWse
abuVarsAqefYAlwmvbam9fF8JWrVqlXg3IhGLkiF4Pgb773qkbKIINSlPH5Tz42UeObmaHrVdsGz
uUS39oJRZ6W8o7eKlZZC9V/Y6mD04m5qoeGXgvjIdBldX/X8cnOCnQm3Cv/+J5BC6Hmk2aOLmIap
d/fxcMpD4W2TuE1iK803vdYZAnfq0y/bc8qCrVbRBmrsf07ONGFL+S+ZShbgmSQ5o7TjX/g22vwm
Ny5EPl0sWdBW/4dkMhzudAL0QkPiyAetXHvfxFK6aDDd5CA/3snU2+OjOQD8lcePI3MdTcdH99+E
XmVdyCD7RuRNipv0HFS9tPcfIq9d3YBIxwT6wF+w9Xd8ZELXQ2aSuOIvOsUUGnw9MKP8CdDhnIqm
B7k2UBMyvsV1aIUQmHtCHwmKY6AlSUUWl9W+lumKH/eYX9gVCEfYsHF0+9w/iLu3NO/2HmMCExUU
fGmZb+FPU/I/X1RC4+OE+QVj9FQMh5CM0d0U3KAW2bFXq1IskM4xpkLEan/TR/FiBtPq6a/5mYb3
XCKQBF+FXoDwFlILgYjwZn3mODq21bCj709zLFYTP6afnB99DZS47j/Tcbf5gkZr9WDr5kzafB2e
omhRCDREhp1OnJFrrZdi38mZigZdPFjqnyRjXsP91wCb8JUeHi8901FhPG9YTCSYvNC5+tuh36Un
knO2lWWiWTyi7WYBH4VSHPElT+bUtGj+umSQLfbamSikCGfBrJBNhFlpVG1uyS89N74MPZtuQIzW
4TVnBnPOW6eqOQOQF/U0Rs6q4NUjcSgkdd5huS8NmlncrbnKHlqN4uM7rmZU4WJklrPMiUTDCzwW
FD9QXUyxdQoZiUioLPXUxggtapx3Gl+cl+BaxL5fG6XSXJGY5ey6Ih8yAY9Ni5T5wt6Ko6bmyh3l
QcPhkeIyFNzHKEO3KEjbK1ui/oVqkq4r1FY1YEWMQXD3rxeswXICtAtIZfIbwgZ1AWV8k5pYbFm4
8C6892q1JMbxIDy6Hv/PySYlxQEJ6u0Xyi1YUWy08AnGBL9Uy8mypTYthN2c/cRw2ptYQRg77Jw9
qeg/JnoBjxLaHHd5/Xl4kB9XH8PCc7Uix5a+5f4aNbJ+29X3TYx57VTY9spMNJU6ShXpR6/7mA2W
nqrF9dR/BYaz/6QSui3b/mBZlGChJNAomwUD9XaoZZ09tfccL+yYzhiRuP8Tt024JWxhlCTT8xNm
T1JNN+R36PF1a3DP6RWgVtv7Mb90Z/VqGi7pw3dS+Mbv7JwlOyWvkdoqECvsISyZ6dMubt2kqAfb
UXh0862eImvyEYu3Qtsd4sgGpBMEpNre96y4fB96lvmh8qjxzX8TfoHtjYuNrLtNLI8Rdr4uPl/x
VkbAeLBdMFPVfsNqeGKDbzYPZyNhjRXIQylC7K7W6HP0nZczQhodpGtcyQEOpXSLO4r2J5b1WM+n
T9wuq3kLlDbqW3ud7hmmr8dbiFa0PCi9S12Ngiphzf/zpEpx5r2hINhymMnsFCkE0Tplyja/u9ME
DZ452AWLTaetyr/FMpg9mzuWTNgAKmGpNR/Fx+Px6O6zki+QKgWmHfII896lMqca19Ml+A081/Ln
c3CgeRdTCA/jcxegFhIBBB1MRRl7VqQnuUMaKj1VO18pfouc/qykgztawIjfmgH3e953vAaETN3B
3SDrC306CnZVmHOYKKbvGozJmhLWt1TJ9K8FCb68fqGO0TJ25GJIk1Q+m+WOLVzY3hpnhu2yPR9X
JdLjDvsP0+O2yuH0MbXGn1EedqidIbhaHVykhl8yle10kFjGLZB/WmsWfmFm/9XmJwLlefjWVXQG
4mykFRHKMOmbCj2ythZaTEu1BWRCZSeQOJcU3kRmntYhESJlZxkxitW8Z56EYVFfAb6n5wY2Kaag
4lyPOB0qhlckq11XXEvzhA+/MSjTOiXL1mPmwW5T8j0nYJZz8D/58wtr1yECuRR8MFZwjlCGTrUI
5sCRknts7R9O4Yfm66DgZfhRx1fXM2pQZwRoHBwC9EVc1gVipnnJupUQHwcRvcQZVUgPJiCO4iEc
YwUC1OJJ8QCSPmrYg2soOGL0rBJQz84pNS0onXrm97I0BLb4vnoaXMaW5i33FQ0W652g6fZ8ob/p
P7fTMSoWRf9mSE28CtW3Q/c9gAikbok0iHhSCxnHhXzadsz0Nzaxk1Bur++ME0TGgHazeNy8Y7Y1
bhZ9oYeWnbzc4SVFnRB/7MKlhxVRVxD1c8xc6RTJqX/nK0pSSB9QHtEBxRzKBJ1FY7d51SMVXQ7Q
o4xA36zC5aE0TAKhb7BC/WecCXh+T9W4xLfla8fcXmsFKh0sN70VXInDL/yL4Gl7h4WuEoloCnoa
KmngEdRDtKp83DgJ8018DfpSbYVN/1XblI/7Ae7ue3yRi4U5KFhl2LMVg8nHQ7UwDS205n9vgRJh
VKWFcbBuKTGoMLzpPzxaCliH7eEzHuT/ocPAWeT8DPKoWRtIYExhaneAtz5bukTKSeSINuUvEEBJ
Vf+JUbWSPdz/GbMSW6gbeZy4Syl0mro/uCd2/NdhIYjO9Mh2D4usSJzVzu3P1epnTa4xK0Gg56Oo
y57wAU54GnDWas4CDmy5RGgnF8Pu7KnQ8NokdOxxJMg9C9C6+FtvzgAX567+XzkDnPGQbXTlGcdP
5iFIGCu/EkVBJjzEPySzrUTfQMlTOpW2aVhI7waK/mudM7hsTdicGSlXyqHGIrY8GJyrhDVJlFz2
mSfpaby5m3DSadQfNXx3B+mXwWRF7wRkWyZZwPrLuC4KoEH4duna+8KBS2hqlIW9+kru6A+mVkr7
o58B6hde741WM0cWKz9jrQDNjEqcfZFC+1WiAUjsG1HOnYsKF7ItWc/bN1TNsyM+6snlOqvzTP/D
k5iOkW6+q+cMhxf5Qxur5QJNBciSkgHy/5fOzmzkwOqXvfsknhUt5a6o1+XSuvpfaW3hSWSG/YG7
0hqaNkmEjYHEHZXG3GK9yw5gILAVnvzcWdxdiPbfRoN03dmxfFenIEWIds5Y5ilThE/OZ6DS713H
TYChlLEg7ZBA9HVSi/PIKh/P2Cda5P60JCZFk5NBP8hrmamKmdc3LubTX6d8jVWQd1tGAvAoDUEK
jI/EPid0LkDT+63fpJAkSFv/SqkwpXm/UrD7HemC195CschVVZD9OZUddO5LtDFC4YblaxqKJLJA
72I1vNB7QyjsCMKjV/KSgHpX/ihjKJskBUIvteVBCNlwseEGAsVeDT1z6/LuOeJCR6U1eKCV0Eko
Tsnx6QR4FVrwDfaLvjiPuoXLpm71tjXzIP93D81DKy/JRncUG2muQAuytZu3cE1qcMmfbD+UILcq
0+yx2hu1rAO5S0tSpgcN5TxtBX7dTfg+YDtRB5xO1lBPXzpfLcTFcJrYbNpYTksrRjacshOQtLCE
sh1qlZn4PG7NitjBGmWGTytggHsApZxghUbtQJd3wz13nFDLiL0N3+wOxPwOd7Ecis8bVdY/gfDT
d/wIDhmbpqgrrF4sBfR2mIWNEYLJ/18mPHmiSseQp7hlZjsHEeGV556G6IxFMvolGRhG2d7/jRc0
KbpGC6t/vi4raU8ZPGfeJUnN1C6WnTHd/UhtC6H8IhxVFnqYvIpt5Ji+Qc1Mu0xP3m1tNYTu4wZD
N2KVMer2vfch7F9ejhdbtml5WDQS7evoSHIwiODoBMRWiHu5SoHZxEIU8nftG1Il6mU7PwNJeUCb
uKdE4+iwqCKqz+3ajemuM/0RmzVIzMxDggrUoIcWQnr2/fADxXoOxnMBRM2SO/a9AmBbPV1PpX8q
WoQJfI2rrEX3IHKUjWa3yYM0UluMF/MC6MCnSQaneCkTZPRazfWonWxHlji/0B+zNI3k1lbcUfdL
2SIazUaLEk7MA/K88JiSqLOSJwnlUBBDOJ5oNJ3K4C6G5t5ZC1kx5Rcz9kOeAVL7jIaCquNQedLO
MzOJfCSWuHTiSgOseRKlHSTiCj/nMkTLM3Fo/rFEKwVlnSXwZgfy243QvGWr4bR73Xu1CbMihVfi
ozy2xFO7H3Kxnp7g6YfgyEmhu2mkZWHa3pMU9G5a5764oURCiO8wmgEzE2Zg111/nzpYdsIO1AB2
W1pv5EZx11QiPe+pDmTWzi+6ipbJof6Ht9uEjKfED3iQxP4Pho8bSDR3D7yPw/ZX557qH/udi1Qw
i3TlBXWKO2SDlxDeetvgxSxgp0Jd5evyAoDj1EjKG6nHXcHQbA4UKI+qH51zcTK0/Vjd78AK4sVg
7g72Q+Vjojm/bLvpS7qiMOtfIC326PRKHUROKGrTholeZRXZ2sopgJT1Be4/Ke6n0QYS5VYektv8
1AzqeNtkV8Pa6UD05DlKAjKCSobXLdTsYGKPvcInJm1SZrhydWkjaSzrB6rYUZGpJeyWBzloTF8/
7ljCoDZKtaYkTCXojcnCNd6e82bBPlJYKKKsTkcCHaCspsyn9bNgTcK//2l/9Ce/gA5IBtxQJp2y
0gI5jf3Hoz3QjCbAO9DkYZnqCNlDePyaboHqTRVLVCL0qqcQwQ4Q+2AM87Du1MmLASwvzoTfJ1n5
yWRT4waQ5m0wF284e6OIG0MzT+pP0Kya50ixnCxk5iYipXM+Rb69oXzoQzJnnSqSsVaCSBtEC5Tj
TyTHMkDH6y6Ez8gmzFYoVDft/XeJMeOOu6NgDLx2lGN7KgqTceSk8pQJLnGYeqby3wbwSV/7ZHJw
PlrO/uiIBEGtsSbJYAw3DkQHDKIBbSum20G91gzhM2GesAHU2jEXPpj42FYKJ9fKDtEmpN/RpQBI
L+7YCyRRciyP4Y3eOI2pmyx/vMDHmZ2M8XrWnu1mPralpNWMJivVD9GExv45ZADga/7udxbkPlDt
u7hpysJ8r44+EosHjNH0V/AGWpOtRXuEHYKS1ZhuTcQK21TIS+OeALdcAU22R11sgGM8G4OL3M9o
zQei5TPuso1eHVzCJUS+7IFAkAXPgUXR59+i6bSTsKh7hz19/YEA0mDYCsNbqKuQ1haxJSdj/siC
KXgEoj87po6TZqR6/DSy9ZoB5nqDK17Ofk7FKoAAcLIZOd5UCe9NEYCrndvfZwM2gyeAvgT9XocM
9bYin5A+bB0Opiyr7YlnP50yOyM+rJpJ9MfRUvLCl9A7cKMk5N9PxYLS08UCVvmWKy5Ou+2/d9Md
T8Luwax2mAInmnk2FcNqQ9LC+JZ57eaki40/OdT+IxgktYpc9L3ByrmuO35MbkOmoUDuCSrzxTkE
PyacuUFN9ptqucXbcz8726wrTobX4kPyVCMMVTqQqlhUsFjkrtH6tGuFlj7g7fVsQJHBt1P5rn9v
ZRzgTGBy8WLRx7dnyGirY/DhXhohfxsfySggZYPoA1dJeMKM6JeerZ4C1Q6TdBAvxZ5Z2Mxdk9IO
5nKH8ZDSTH1d0QH597Q/2B4KbLPqkrwxcxt/15Hp/HAyFAbLIgFcZq7qdxQL+LiKrOf03TQkuQdW
T1pgkL3PbZiIXYlZktgQfE3CdbdKJ81IPnWqOZRBmoxIMyT6nOAXHzk78FgieEEQ7JgZ91KDUh3Z
byko2ZbC4nZ1W6BGAcQDjHFcRkhTv5GKxjvMZfjabBaHY9j0pm3m+oCTYCTO3zPcvsMKhi2GaaMW
/63f1C09krwoTPpcVdLnrX6TWOtUr9jHfAtVTYC0mea0VVNxNxZSLtHeNDq4kwH47cjHvaIiV3NT
VMKZdqwv7DbhARS3MChR9sK6Rr5zu3b5HCTobFuvrnIfUXCpPw1oy48od3k8drlxFzBGzmd+QzN6
2QQqiPVVIA975L6RStvyTZpc+W6Ik27BH3TjMf2vqVHDZHjEBLnXG8cek6frkMXPsaYCuU/a3Y/L
bOtHfG4RJ3Sgk7dfsQ/Vp7/H2SxevGg01IWgr48dFlUsD7GmSQeD9NU2E7mUdPSEhm7yM2fAKKhc
Um2o38AceY0QM09weoru+gMC49kiqgyDFn/xikgZNXynpjuHkv08jnUJKbQ58Qso3I1XljzJxRF6
EGHZudWZ5mIJOYR4l7tYpvsh23jz6mAYI2XwSJ9ODIuSlqWwwg3CBiikkK5zhtpYlacOlUJODXXG
c+EWIVZtSiuh0aj9oYZP/f2jDPrDe8iZAF2zpSQbKkh5ePdxt1ZxwulA6ztMJwwmKWVhw4yErm8j
BTnvKK/Rv+yY1yIf+tf69N+rBIGxB8kOPx0FcN3oyZVYDXbp/S+kmG7XGxuiqlzRGbgj8klTozki
C9g0sKhlpI7jSm7w5yGs1sOUEGbB5ig8VNX15+z0GhC86XEITogF1lyo4NSXxNx7Jgt0FrGDB3db
8HeS2fQ3yyX1cdfmfMU59eE0I1olRF7r+l8Rydv8wUDXFwndvRRzhkM/bQbpr0ZXAYNAS4dJ1oYU
vv7oBxjKB+mymqIkQsXkCkjq8Vndgts+bAFbri4kyBKXkpH032Yubfz7d/oGYrpuTev5WxjqM0aA
89rYdvd9uduR0R2qCssDycPfVffQX108ig1K/GENcYL+C7iVjr8ZOoY/QKBe44F3fPxW/edQ40K+
DKOYIVPREZnplrmnJ5jWMMK59lwHvkxpdZ9QC7+Uyxt6gb2B+sexNSiVa2cA53Au2RIugrRcChs7
tPraw7u6/g0ozTOWVvXNdaUA+8816eqViN0sLV043Al4RjSjAORoBuf1Jn3UVLfGHTeWT+Q7rAN9
crINJxmgiqjkB66u34v2JNbUc9IsSieVWiRdShfPCdAv+ArgKgD59pWhZfhpXKHkeUeSBQtfeAXv
wlecbXRAdotkobKtMeRFIR4MDx/Ujg889rZDAW09qnb8UBGeD7aYv1lThupP42fmcYzLw3s9I8U1
Y5lsC8FdGdd6Jz8Z3sz9As6+8ICpr60MzPa0r5oypQx5BRCeeRex9vaXOEAMp7Iqge0UTqBHe1X8
ldeSnZGLRJcFsL6XPj+Yau/Q9CYbiubUtBByqOMOwsNjpZsqXmbsa6oZQA55kpzr6Ae6frSbokIU
3siIFY76QTmlC89XX77vmBcT7+LNOYtoF6izy74+GSslG6kljRBqlYBWHRsOlRiQ7NztRXNk4U7i
ZaIcpZ91/mUpx4Lmugi/pfxXwB7I7uHt8BRd+TyZI8HpwMSFgrlU8Jbrbpe70Lh9aW1j4uDT09/W
W8yQD9FTwQUVvry3e5rR9ocqK4BR/39g0Ffhy5ip9iVYNvki7WQIt7gWjl29lnia9Drqmd9eA9Tb
bD7UQkH/VXRE2E8zl9NEI/5QgnzYpE3OGHxBCoON8YVULQ4bwlyrSrzcq/WwCgccpPBTDuKnkIZl
BfSY7QoTGWDHmmaFiKmfIkdzHZogYmsxcBgieROgk121uhpb8/ZwT//E+eYCAgr+tnP+0IjfKjyh
OatNsmuRpoJo4YnOnDhSHb4TAZb7EkpGW8eZgRyXkoMhqLMvIPCwMuMAYMgRvtdjxZxpRj6Gd5UC
VTYP3572jlVLOqMC+tPmLDENKAeOn/gg4t/tChh3RpulIucaXJ4E/fPea0kPtADRyJPY27Jg4Eyz
paKBnvBAU62CZJrXhMIvVNtpy9Vj2dR7k928PIRq0zTtJah9mn4okBY+NHcmD+avi1nrssijrH78
CflesFLGwrYQSCqTFWX6TZxu60MfbltIL02yOQdSKV7bQEKxNIsoRjjENQjMIxLuDdF6LRNxwknO
XASx4IT2PSj2zNuh6c5NcmoicnwA/6QzESKOakgrKiCPu/p6VTrKHnSlGtRFX0UtAeHwYorG1bW7
Yybm2TNChdESnFvoPgnanfts/Rt98kknjqx5BzU2qmLNj2f2o/IAk+HnkLbTyG3h/pAg6a+ByZvB
h7bYzpgbUIa0nzs8hwRdf5L+wTvcLodryiVM5yGQ/SX4BYIYUmPN9HP+JjG3VSY1tkFjPdPA2uqn
EnXJcjKpi9/ydnWpsWQ2G/UXZdTFeaQW+SSQ3uHgn5tVOe0aqLHBDSVSha6g+Kn08qMKITWi+Pdi
g5x4wD9FOzhjqHmU4ESdLe7AkLxUXHHOa4yAGafAbV9YpVkOzdI23zEN+rf31KBK+j8eftdiBivu
+yLqbPPwCVU6jP8pd425CpKdN/ZNuduNIUOWqnajJdliN0RPA13nlNaK1XGPLvszWDK1yJgMasRa
YG2MMRvFi5zl4JzsmCQVjm0744o1mdfpkeGZL+zQlhj6oAaVtOaytlQ5VgQpE4qdA2Z01/vIbH7i
FUAt7qDSa+L82lK4bYVqjpELzoiV1QfBSQxhXAIqgSFrLL9McCC69XPtIp5zpxfnaW2W9GUrZ5s6
i2PrtWUbT6U/Bp3oC6dSZeerTJmUEYC+yyaQrJc2ZKl06SNo60QdzHqTyb94P2nG9xWoIIcrU8jH
6ZS4npWdCdJ5EZ0hWYitlJUnwGnYRfMiImWeftQpxMrVlkGO6e6LSuSqP+70GkPr8GtkhFb0sCEH
X2mlmc+347mXHX1Ukg7Gzd3HvEGXmqa0MDtfHZ4Fml0d9ROBsWv+ihgsOPqyBm/KDtQafhAI21rL
Q3JMbbDguxCY7ugb3iWBqfqy3RBqGr0qidmXhsuVIWpv/1EUe5G+65i3s92/E/3zWtKgaX2M4l0T
o1If6lgHAP9iTD1038E98IQT4jHYhGBayWXYX67nrGQxTMqa09vafYGp41aFvIvwiNMMm7DL4x/q
nliNiuQjmZ/r8j2FyzNPAtCUPLzlwouMW/fH2B1dEMmhXf3xngBQtN8judWozKJIVRfZ/xS7i78E
OjyyYn39oQ/YKdJeogk9qwIWvIs6VJUPsTvxr98pnctEPWiJ2YRx08YWpc9s92fExQhkp5XRg9jc
EQOXnGuGU6SWfP7R8TN3vgjPHpBe5E2lV6J54VuWfyLWF07Szvm6rggoY/LtdrF0odKjcwxQN1AA
e/QG9jXwtqTyJ9Ph6xIfLf07M7xlt2z2/cUaeopYs4YiCEQcjGU+ptOzCCcwTTX6I02QvgT2r2Hi
tYWgUasMRRe2h8l+VvuI/0wHVkbE1I0DDPnnCVo88j6hHg2k6Zu4DWSk5zDFZoke9bUdV6WhqE8N
xYNQkEIisw2RxoK2zAqywZ9JgfUF7U1Fzc4YEFylvNlezlOf9gIuA4vWBmtlLck4+w90LocUHjsK
Os3w2Zv6dU60i8zohZhVmN85lhTuwE6MqNEycYesNHBKsoN17VZ1RCw6/beQ4aDh41VVgQhR9adB
0TOVX7HjTzXwG7bVD391V8aZooLoSxvv2KDvbeODbbBmxPSu4zh/t6JdyOGWGZOyNMcmZD5DI4zl
zwQQph3gqoOvW3lp71Wlv6s2h/H7EOpvm/86TF6b6jBt8Yp2GJjqK+k/vjbAv9/zi7jFmtcr/Kgt
JcxgNl9qsSk3J0w7oq9gflnbUZuyQxcqTkXbtEslK/CaYXHpMmvLcOPOOhH6i+1jCnWKICGQSANB
OYSLj7wpJ9eGvxmJsHXyyIy+V46dMTyblYQ4KJOsKQzOgqpd3ChSu0mfrir1qwyep1WtgZdZ/JlP
HyZP5oajqIuS+CQYHRszSSVMWkDxVOLmfLHuk23vSYimXimJ8Vo0joPX9nHfzZFKk/YbQDgt41x4
hBy4/V5D28kEHoZvd+B+pScjDfG51Yw+YyE65qTUHasiEJZDhwE7p4oRJCYpvchlC00JAdUM51zR
kL1f5894nQKW909tcdb7lqf2J2GqlUAEKq9+4jD/mf6MRz4zUsgFhMFO/rwU050DZ0pQVLr+bVMN
Nu6fqv4kWzedr5k9ZrMwy/PryipKp7vfgWQheJNkCYKsbwC02EBcVNVC25aWolPbdQpD8lg9I6uT
pHFgkqEmIMtOGT5niLtxCl1xksTXrbSy4QAT0/aAxCQujHMUm1wahADRb31sA/HFt4vASl9pFWnr
nhUwmlWg1RC2VaErlpBhbe+C4ZgN+/pAuu+zv0dZhqmimzgYgZpMoD59tim11Eh2y6S+SN4wpWen
PtkRWKKYZb1ghQZ1lbx2po3LIOil3xqXeJMPYynFzxVMmrBK5RLki8xwEx6RZqrC4yDbV9in4YYb
JJ6/43p1VDC5zaRbyEZZR12FmSq2IvGtdEp7GVG+0nKR4P465lSFUsBYPZ/IzIxAW4LBNnbigVtS
SRnLKl2VefunWaQlwa3Qy3PmgA8FRyxv5Ol6thImS39dHMZHigdAyxzD8OamhYZlLPeD30/x0/J9
wT5q+jLjWCDrHBvZrYsoQReyKM4wOFtHJ9Us076/7DSLxZXgXO551mGNwuYquVqe4JXf4kmLKPQN
0+GVe7vIVWPgTp1pruaKCrbDE5c8W88hxHfL0l2E2l7/Ds1XQIv3ApMZicWWC/k9AqONAoFW7KDb
tCIu72wELr+4zrTQDjjSBGxFw9+vidv8xQFUH7rGFXxWbP6GeHCj35T1zwYAux6qN0mmcDxGp0SG
omafBRNSPJIqT4+DHoS478XmCR2qk0iA/Ar9CQuhexxfOiZZIiIJfryu1Pf1sm87C5bPGYfk+qdU
ntcyIv696QOhPyXOibgFxN1dH6YqFNNNL4Jx5CDWKdsRNlMhDSDvfmghvS1InM5kETszWQ1uRfWY
clTbq66riod/WHJdC3IOUzcHMOFnIw3Xhn8cb81MQLgJQZBqL/3ZUJeAcnYQMMRoxSSriBsbvE6m
hb7DiPHXV7hVy8A4Gvnsy1IZVnIWUaZF2mleIZFwSZnn+VZsjTK0wtatGylA9N5VqK9EXAFshIyC
Ox13aFKlBwqwDhK+bP8cnGwoCp0xZcZFv5vL39FTiz+9UOUyt24C483jPMVan3rrVuVQLEQB/O9I
tkuLzxcH3ceNnDcNmrhwC+Nc10e9V3ayNDutWdvphSzu7ltp6BNWK8/YxSdPEDCbM7s7Dv1AMybM
qix6pAHvs22itGquH59JHt1Q/snDT361+UX8YYOBMRrIAMqjDPYWe4sPK1i6N8+IOe9dwdSkFpil
F3BywxXllnJ4YApz8SBoiV0s12M85CTs/foqNsS6Yt/1UeHyYVzTqFiOc0utL+Shq7B5nXTxRmde
rD+9gsQftt1LhvtPcJokkG/2H8LORQgoGm7EIKivrBpcYevINyViPYkFiTy1vgBpqCEKSD2ie0Sh
hOFbPuri8TBq9ui5wQHkJIn/VMvxs34ZIHlMLDIskjbIrAX1fmcc8v7CL5IFR7wL8RS2HBmXrEQj
L39JYunNCNDqc7I29zmc7TPKUSHtdld9CFph0icoC+7Akt1tIOC0TSlLKn7CmoXhnNQELFNUhlaQ
0NKDIUu4Cc7V0mBhim8+BxSKQBtzapCwU26Ojcvu1J+4lryd2z6lTo5wadI5o79uvQ576vy4F0Vo
i3ppcdpCTEmu41xNmLGn81XBaWmXIrlcnaicuVTl9JnmOeHxWr+IVKS/v/fPjh1Y5Zm9+XCgnsZe
ervvBbr7HjpjnIQ654Na2A8jqChIcxUVfB980aS5lY7A5VO8RpJsjI+JVvtVKPnRPHnQ6gtEtksr
rKyRjcghhRGVUtEz9nNA6kYQ7i/fQbHALA4TaBTpBsTkLJJ5M6TVwtju1jbwyHKEZauGGc6wvfYI
Rq9vX5O4sCv2lEuLrdJeKeJS9f006xRqmXGdWjKbKJqgGQcL/NS7kCghGVUIJHj7WSxabSA2IiX2
QJxXain+HOL93hk6NgxJElLfbuHveTja6zdP/Qvik4ABDFLFOhRvJP1ekIWPkkXG95VfMyDPZuc/
eEpCOGYZG11CB3ecBeCN7913ZTLBSyCIdGmtnC1a+9nfonfqawnG7U4xs/bj8TWuRlaMwzzjvACK
Sv4/5F1054dM36Ta3w3TkClnjgjkk8EK4bFRkdwjr1aczZHcYZoO6YjGYxeYsfVV4tyhyzOFBnKc
ezpcpY850lieWFJvpbXaYzpDnKOs2FFLCoqenXwU7nb9JcWFTsUppFImSCfM3AdgfewCb4HsSWRp
U2+Ls9LKkjhp8/l0XhQ6sW2YD/0SC1lDW6NYOahSpoqB3eYb6OY4gZ+5M7lfsMKxWjjsNdn80EPD
j037w+6HZfpPIvWHst7ymK5q45XqBJKkDIXW+Cg47UUaOEaWryuZ6Yg40CyK+hOhi9aCNzp3eDEt
CJP9AYoyZ0Cz9P9NxZ+Tlr3BSnh6yfB9ZY7RFSvVhb+dupwBW0RhN8UIqeUYo+27h+WDO99rNjUW
cwm6W5MMBlii5Q4fUrMSbkRgfF2w1r710R20h/eZgO/1X4z2vpvp4gU+IqA2oy+eg2Er+pNX6fKz
4/yeMg0+5mm4g/gRBfaaJxLtgQ89Q7tWP+axvK6mqZCq+aek07FViFxh4ZyR/HLqbE3RqMm5Ha2P
DVmulXcLEpFaui+DH5f+SEg34ZNX8l+ztH4cyxv1aUbzEapYaCLMNbgY5opFC9p2vMaXyGHKE9eV
QtzjrBIUEhPl7QkIU/EBId+kfrt6dOmzWVk1mAmyHnqyiKV2125QWT6CAwVmEfNw4epUSuk/2hQN
a3L91LipLin7avtFUWZwvaeW2jgIciFUZswDcT+imrIiGity0cCITcFWbluG592PYOcUTCj3MYqD
OsbbvNVr/HW/mg2R4AI1UdyG9u3btAGn381niR/F0k7RwJm8mBVoY8lHJeSXIQUd11kgLqw/NTSH
7S3UmUv06FsZ8066CFqMGHllzTQSea7Gv/12VsnxfOV7KuGmdguqkLfFarw+TLfz+6gA+OneVWAa
KEnRqMPJxCyzKqyH7d2BzwT9CRolglyD88HDaX8vZrHxSrCSkVfOG7OgbNDmGuAEevxGFjZ1JVSn
/yM81tU6ota5KCAolQdTaeovVDJEbEhwodxFp4nM55WWn8+4Mvz8lnN8VH1FRIlWE7Vfa/6vLrT/
YE0axINgWZrlofAlEXTae3ME37FxJz3xapMrUd2PQgmUA4o+a1aFOMuy+1J/J7h2WSleOmDY+nOa
X2Y/6+TsBTy7iIm/P5AeCwGdYP6GPssVpoqKgS+nwDy6CnSUgCgLxXCaSm8Jsn81gRBXq4jbk346
v5G1zRNgR/7CmTC/CHFiDAj69fcTMwt455xawYXTAEwncxmb9Cu7qh3wfIcuDShtF6oNn0k02lWT
CnR7sPCbMXCQ5QUhe5bBqEloYbUVbnDea4sdMg01So8OW8MK64hAZr38p8d5TRk+D/YdTMo8h1jS
llF8U2iUJ5lOiSh/jCoYC4du129QEouwP6IpXHeCQIx+JupHTaBFammcAKy54RHjIFz+TPMrsRFb
B6VebCCms3wwfCiICvPVZz6EYggUefLk4n5RYAls25iEzxtG6AJIOS0ApQlqzN8puydx7t6d8JYw
OYc9gHyldBhJ4U7DAEzYJtlm5NuTY4wwfXMd5VUIIGSmXlAoKRZn/ofxxzSJeX7y2ZoTdb6gIFxB
qeXJikFWvBhehU14/ea+dfjGoeGpsPc/8cuRUErDPhSqi2kvhqS5cXLdixchJJeMVI+dXVTWNEwx
umHJxBvUCaxUpIMwtTJydcU7CWuL6LwrXaRQMVZa+r5JH18JqUEYcltkKbhvhdY/KS8y1WDpMLif
fkXagUmJ77PZjCktXhZyTy/1RzhsSSDzE1zsdFbJRukN2a9JlJdJgtVQWBYyApfOBivzi6dJVN49
e1wy3M65TpYg4uz+FqnVZcdXU7Pd80My5xydIWmMGb3vhXYruOyv9G4jFhfxtCUGUtCmCeZfm+Zt
7WqhIP2UAKoBKns0SI5DsypkyaDMU0MVOv2XNBpMsQYJ1fOFeLOO+eoZSbOmikeiFYNjYLbmLQHW
LsYZAFjTAeucOn5bQhBPIiWxIDE+07tki+d+b+6EliTcIw/H9jHwDdkswCpZlJZOAsr253Sl4r8V
bYvE2yP+aVL2hTbNdIk79AexM4SVDMRLo7hYoSjiYjVdJ0cchrK1befi5csYH4pNYLCObdgdYE1v
C7jaJrdMckyic96bo5sOssPPB+qbVzWVXCTEUO8AlF3Rj9qFo0xN2tTCcpZtHElJ9nvHn6gtDUps
mqDipDdv54BHaJcSpwBYpxPeJ1cz+SzVY+RmJ1M846SnQi7FpFAtkjgBXfu7lHZjDu/7cn/AHEp9
aCnekObJdot2Ucn/Jg678uhnbFDEuNXha9KjtGPFErPvVoXrSsZmRYClyW2ElV8k0/IXIaa8Ll5S
jSvMEMo+3LVN0a1cOfC+K61WLoZXTA0YUFu65HgmcCxexyXJsIBRsNQUt2+/7GC6gREVqpbwxAC9
njI3R85wEWYKY+EkyCoFuDd7I1gIpGB5WzslAcu6OGhtlyx5uqzDUQxUctho39Cg0stB6qzJP2AQ
vU83SWVll0+GRNVoSFJQ6pl3HuyMbofz29FiUczotNG5XeW7VsNETDFzVIRSz7bq6AirvXQwJDQ+
zWUTp0EgqROPmo0LSo3m4weWFkZ4vxLGv0jjRVPPe9vvedSFSXGjhcBWC+Ukdece9kD0bzstg/bP
pk374Hxd2gZ72DyF99pkS9Amz5gp7WriqmJMTvU8wKOvOpu4ta88WycpFthdcNZUIuGvXgtUgTpd
fBNiTEtf+KRtvTVTzumBIdXSl77dzfs8CHZDqT6C6xhU0yXCNMSWSI+HbZEOZPBz3+rJaBpbXGpX
UpU9IWaTupD6KoLlkdX7O8bdHIfxD9SWVLOGQmzVTLsSph4YNu1f3fF2ucJ09Lsr2qU2GCK0KzOP
mEORU3UKnoOcWv+9VK7aSlEEcAeLYCb96qWa+0KBSLW8D0eOioWHCQadu6QE2Rkhvu/QWMnZQBim
hRH5gwFAoQkL0Ru9BudHIg1//L0fu4w8fj3w3YYbmBMnckTGLLRDYYwQtnCeNwLsqg+IigSPqNXS
o8LP7ctH5vF3NVPxg34gyRq7mGSE7HerSsVqCWL5kgKRjyjI/EknEWe0s/YzdOKf4fNusYNru3h4
WCkceJMZSpyJjtipVxeDcq2aBt5DrG6a4JwZmVQKvr9kTXA2TAY6Wi/q0VMmSTdLo3BBpJQ5Gm0Z
2pLkeezuN/j8GaSnAd/MjfLos32QQoVzr1DXYQBCvPKZBMpwGEsdCGQauGLMo1pqixmHDuzqp3ky
iGMp1gX8hcmrOHumohhWX4LlxLCDYgtJ4V/ftjBkBbhc3jFXub3xXEFbW2LraXkRfla7KCluni9/
C2noEYqTKuHIP16Lu8UfTT4TvMh8rce0Nri2MpYtxiI+foUEzHO5zDFcniOA6rtvfDqHEz3ogV0K
id9epEZLr0cqz6DwiyCjCilZh06WopLx+e140MOocF+dFDOK4naWUASMU78M+HJqm5ZZJUju8izH
xk7i5R+B0KSS/JN6RcE54b4hjKU0Kz20X/btDy7GGNHz4wGK/r3RC5K+LOg/1FC7335h1dsMfuKp
5Oq8ZIVsjThNCBuzEvnuIh+bzq9dc6LWqE5hio2m4BhlidZJNnrp2Xv5Pnq8FnCEvgVP3dxb5AnZ
812+fIs/vBXTpsT2nhNQce3JJ2m1bQLSg7rAMEMfp67va8vztT4Tub5+EXbNKTLVT4LKnzLCm3DL
t8xggn8EdNXu9g9gZffMtnotI11kbQs0xZT/TcYndhP5rzcy08rjYMaD/Qi2TW1dWbZTEOat6XW3
72ndQTsVgjTHdQku/HUHAOvu4jpJxT/AF4qE74P0ebW5UCYA5VAAPL4vtAGOZ2QGgCKdSebWunla
ikVrBEi8eYXoKEn4hW2eF/gaJxsv8CHOgmw7+BiThupN40ZFSyv1kGOkTPLgY9gSe1vVCdvlNkW+
bZPXgubQT5qXy5v96+hJ/RTedh21ATyj9+wCTGvcF/GqY7Y3KOa+mntABHtlqKescn0VqmvwZF5r
syJ+JmqANH8sGgKiNGxmFZ3RJ5r66L8tjdi1uJLKnMA1J618BCq1k+vPzijV8SOSy75G1CwnsY4+
uF5Xud8EjeAvp08R+aHe7XAFQxn2DN083+FTcrGYPyYmerH/KNmbFkiswHZt3zi+kiKOGEWIitaS
KVe/rLEpda3hcx7oVTIBJL92pxAzl+vJbgpcE+4sOArzlHhfQSTFmFc8Jjrx8u9aQFPjUiYMORmV
RkRmgCnJaOIKB8RsngoArsoNWwGY0LDjMi162xhediursL0It50ikoVUYkfwE0WqoA404llrhqmf
R0KKDig9btYJyZYnXQCFMrW1L1qtc2dJZBYOIcgAjXi4R/j4jha8sckorl7uTTG4XeZusJdqqQxH
EAQVDr12ZUTXaUp7nsdgpZtP1itaVvGm7rrFFwfQ3Gpa50+Fz5N78BXhFdCPRWDww21hUgSvWYsB
lFuHjBmkChHvh2dzbCmMZn3QlbgxTP0bsIoy4koVsWBi9YQAzvzEd5QSzHHN0QD1/1hVOYW2ghCi
AOpgppo5B3XI0MfND+zLBJl3E9BLHy4V79pO67LqQGLIumYxMbqxc6CBhT9e8PXWfDQVykXlM26m
8Y1r86qfrJRmuFrW0wt6p51DvTnyBVH/0chxXVltPYypSpRpZA0wfTR8dEncFBmscCUEMPMV96Ni
CZkmMuI0YlickKxB7GvnXEpHaOIoE2xLeuarmLFD9mN1X9ECRzN+GJtNqyQ/NyRhH0e8rPBBrws8
YKonsZXxPMtLvVqI2BWdJF2yqUplxOJKgQ/dl1oUBuG8XyFYfyh+i5clbr+0TvEDCMZheBd6pLbe
3Mg/QXFs1Np1GIUcT+A7szi5VBb+60qHubN+ysoNy9j5f0aLDrmv9MxmrmkSfwuWo/zGB25xdcMt
bj1guv2023y4T1jn6LX/U3P0C/niU/uuj0+6m7zrXUdr0BVyIACDbsGFvMyYEqGRm4RbikBDj5R2
/6qeSXlJgBG1OzIbEJA8LhhTpr/CMQ+WrUXhNab2J0PzdvfeBqjKZMSonVnplmfWTt02ljhylKYX
ZtCFGTf5EBIEmlohE0TsUl+6Pq73VL87jGZ2j5BkxQ9nkeXWhz75alzj6QqVsWqrVBKFqZL2prVb
DQEio4OD0S0OjGdlETkvud9SoHdpr2ZEt+iP6C0e8PrpFEuxdSldmjflXrZg7jvBw/6S87p9nh6F
fIQziq+F3uUldUldpqLtmuRdzyQCnFr3rP9gE421rUzbaab43hpy7S3nhIaxjy3ls4qnmQGbjJuU
LrHNp+VJwqv6N58LS5jH/N1gUovY4KHPw6aahM/UWapgpoIV5tL7S/BiQxaIzN2mj8oGw4i0eIUp
iJr8DjA5iBy2TWWVkIau/vkZE3CuNc+t5yMNOhFQoyspILvdJhG1yqCxhLELSpnQ2lTXFz7q09vN
m2nof7gU4zGpPBlKD0JCRxiTZ1yMv/ljaWcvV+THAcLbE7wnuFInkNTBQbuk89T5+5ZJeGW7MZHt
B+OItY9fuEy+SkZ9ekssr51S88n3KOp8hFeAflAkcQt4c+8WWv4eso1FFxbfAlPsaBNhyzYsOSoi
1PjOvSHq/1wXpwcEyRMfc3L5D8lB3Zda4x+PdcvW4tTT13sqLk5HSY6KaifEpAFHQMrWzaiKSh4i
szrjxWR4Ze57WdQvzsjnCvR9ofn7ZH6HHMJBlqRQx51ANa3Hveu3ccAk1POUPGe+jpN/5/CCA8WF
s8aQ9uhb/sG1p9gaOKeVIt6JNKQIgMwKjJatMaBa3mWl0JrYOl+8N0fXJvgWMD1ogTvSF8ZVBJTw
M7WTGofeqwpXZURU/BqtcxYjQwK/0+e/xkTLMY9ktC9aBPFDNQsrWbUi8qyWA52iUlfy8zNpQ809
O1Q5ahrYdzrzLYsV/rR/daaXgtELTbJIedUw0o8HFy0j/vWJ5cVkm2P4gEqf6Pyenr5rnhQ7aiVd
hj3fY+NYu+X/eVN/h9FXq6bP72t/tF6QuO8CRDt5B51cu/gox7jOUkETBeGrco+KM18fw7Tg2lte
98l2K6RxPTPv/n5N4bo3L9T6oXoKvLlWF5PFavWL/PKajUDKSMpi7d9AIfOf9eIA6s3EM6WwTvWk
ecONM/84wnkI9kHEOMKzheiyHk+mMzOyZNIETKkY4Ip/GVJGMS0inDL4VDQRLBUdCqSOiBMMHd4S
MwCIm1e2NwlyvSqQkWFlLxL5xV79XbmsYSi1bWkjdZx82YU53Nx4XXxU3iG18zi83RLBZbndpip9
j/5kICnh+5OugZw7EdnCMclBBjvWZmF+AFXjdnhPVBIRRVF5CJJhZootdI2lFTO+q1GPXtSkQ4jR
KqW3gRtHshXI4gVrKZWzVEx4g+ZavHyTobMbBhZE4EYNd6MLK+kasybFwE1gNQUIvqySTOzTx46l
5YtjtghKShyU0AMO3gK0D1CssOPXsis48TwHp1pcTJyDSsWwtEOcmxpyNXUQNW1SBqKbShjRTbDT
p8VFe51+JvFA5Pw146DlEmdRGAE0FjZ61k+CuBQxEDcMWFL/KcYOFPQ2U+xPcdKuCKeWOYMWaTPW
onEqXfp1Y/JPRAq5LVWATORfUa0duFR6VP2TV6yaZf7lAJ3qh+f4mFvTjuOempwRnPz9dGWVLenY
662pdXwaBe/We5j96FY8wUHB7Lqdf9yyHbh0d+FLxxBZsWkHzScl26jWQh9CHNzUwqUz5SB0FILL
qv/7XZ9pxJQEjcRxLMb1arjgLgtZoTOz7oDvghsJ1Q9ZZ54AE38DTxYwZ8SHkLAfjqPeH8EwQwSk
lW3bbGenou8qKT9tgJAYtzRFph/2v6qKozhq6N6Ne1Xztl5+N3+mZvV2+dr8JOQSGEb0DXXw4Mg9
4NFbi/BeV8j5GEjCmOrMGBYkulKyjW6/Ova1ITKOOMbrXqjafQ8yPRI7B1ie0+a40+oBg8DClorz
t82JpQoTlmsCFgi6OBaNXMNcl5xtNHPOk/V5871X8GpNPq2bv4YvKKk+D5EjDPXeUDNZQ499khfp
A3pdQDP5NZ4dVMjPznctLKzIGosdjV5TCy5CMTz4ASyK/iuadyJmNeO7jc8fc3PmHwDtk6JQU8pb
03Qjo2WJWwo/U4A9I9UD3qXM2IdJhYLkCPywslVCJ5aSHywcmuCyEPUgeUl0xzn67uHbx9d8dlSu
MvgQva07tsVksHFqoNj7BhHN6H2TSBwMB5Y9ugx3iTJFgfOdezGuFzLSgrSosjoOKMTYEL+4OiNU
pvKb4bqLuOCBxzDs3vk66yog5IZ6IgOVJWXGmvoSXlrnXMT3HaPG+ZcQUnZ0bXUgQlcPjUOQxHM3
faw60xKleZtKmbA1fMOet/xjEexkMPTqxTkcU11NGYic+tVQ44ZB2O9/GXrXZfpBwgnJ8Vzf4hQT
YLnbWm3axEpG6QmQMh4TQ9rmNwbrjVxlXv/x7YCpxN+npdOSUHmT3vlLSgDHc1TQRsZJ1i2vvJpw
l1nfkXp21mkjs96uiIuda2kYyMg5Ua3Cs5W0M1eaB6b/9CNgNrO0Jihfp0cnNSZf6Vt9zgvzL1y7
uTG46p7crX+zoG15KO0PiIDzr8jE8IEA1Kqel9ouw4tbsYrWLNAo9ldIIq4u4LqNq8LRAiH8/qxN
g1nffTz9b2cTFTdz1TyHpIZ7h9SWHeK5NGwmnw2iVZ1h9h6sY/TFY6F4FK1K24pPNSN6bfa9TkuG
nuCzqrkyRqMetm6bP+GvbQf2BMGCGGKrY9yQE6OmiUXl0oZeeGjs+LTlR2GAR55R6/5PlTgRnrMv
jx9eQSfcaB86Aa3Orn4cr6+PjokkDHwu24i1n5jxCP43XBDN98iJAYcIvOAIaWAIK5xNR7v5kJqr
5DSaLghwjRwRDtsYE7LEVitiEZMS2e2CBDOEJ46vLHpJ3/wFdKJpQxo+gmyrueMfBKh7EO4PJx9r
isETtpXsg25vOfM0K0AyLgakq883tg0hEA6YQt9uNibJcMNyaCnfD84846s7L90tLGmYF4pZy0nX
Yqt689s9sdKwwk5Tt68Mn3XOiJegNFfuGrNnmXB5jgi8vRTHmnuXTMSuRDx4OWT/hUGBIBQgdaMH
Msp2q3M9bqodJ7Df8sHDDOnXqMXqyVOowTsdX1C8qt0CKgNp8q1d8egOE2EayXFZnfltWF4MqBK+
Lm/UFzSPtkTk7v3zZMLzHqCltcBTK33OMDWotqfKf5FHyk3yIZvsXC7SFz6s/Srlsu6LOKLFVavV
iEkv5bNJmoGA51xeJSvinTEu3ssC9OkVjxwz6sOJjuMUzn5bUeAUdqny6sP4zpFBGwCRFEKk4Nqg
PddHSfd3Gt8BV9zRghI6NIsyGG6KiknXi4pYq8lydk7rzKx13w3jRjddvkxvFq8XJCYONGcCoEhS
+aDMwr4Rj/bpq7hxe/dyzFwCqsLGxJrWFYdQ7dy3sU35pJbO7DOCF4JRDh9h+wuZBVzt4dikm7ze
wpyKxl1hykfK7lIrA0gyOuFKFtmjpX4nSD5d9srdhgW8ztYBuhn+mCo4JuDcJXhRML5i93npGMp8
vuhKqUSIr9hbM0fwyiRvQEC+X+Y7kLQ5ooBFuAxprGXFoHb94+9PvgyQLD4dUTU262DpVhpeW9ts
GtPW2HQKsR90WH+f9RVkL03k+dT6bIMyvcCPchyMuiOnrtk0dJhCK6Xwolt0EDw2i+lU6/xOXPZ/
iy7rQM6v8fqO8GwJHHAKQnwVSzcuPla+9OaMsLZyEk5OL+Xe7fKGfcdy0buqa0OwpUiQO09yaG2c
KCFS6lRsfjV4SuyjBJ4+169fbaTIsDqvlaEeNs0NrUjmwc6mYhE2zy8zR/eAHsXOFgOuitCKyyZP
6PYGYR31byhJUsQPC93fUzPEZZLVvMCtKqy7dZ1+nQm22uEZ2HTEQz3NPK0BAQ7AK24Hcoyzeb4K
u6hbhMuMdE/UNtI7CtV6KHCcKb6vabLt5w+S36c+a7Wys/Uy2mo7Y5NbQDYNgZ8tPncACgXIubkX
S4QTlnbp/A3IfT7YqlKPW7M43PqphtgY8UOx56dmSpqKslAkCm044yf6B3Q0gxFEiUGvWeofSrmG
nBOxMa3jrg40fzkmWjNiufCBoQx/9tp8d3RNzUZ4zc2mBI2qlkcpwJwZx5ahf2IaKOKJxqhCybrf
i062v+QWnpBa5ieMT6/SIoQfirdRmOmCkztEs4PNj/nLOnclIpBgZZ4vWRpovHhS7QeXLhCjRXM9
9G9DtsvPw5qti9JQlI2Nop+Yls4xWiO4EqZLQUm4C14fcwG963q4s8Vfr4FnLGaxbUprytA8poWJ
tJ2x8SdsDqYE2bNJrvfTD7H1kjy2ggZ8EUH1B4YuuZCZc1yaZkF6n4zzcTDZJSFvXYp6a/yjdqQD
613Meysh1rdTcah96DaYAMiM6cYWRMOyT0CXVowtxC9VSF6eurEqbbo/d4orsXtBrdAZesf0m9GL
RR75sHXY6yDDvOIUbMJpYzTbCnGPMbNw633ISarRbnXOwV11emELh1VKjAQdPXIFhbmZ/VETvYID
c2rA4PvIbI/UP7BrE8GJmSDlc4E5mAm9pNB4qlDp1MJTg4B8wIQX7PHDqdeIhn4E8rBLe69ECPIz
o79uFocgcOgyWBxCjY59Bsb/wUubeOr/gm3Ey1mIEVcZQN8N61+6/jgsyOmwIumbGjFeSptueoik
z2YxbXS5L+a7j3v+PtufRbA9NqdEzwnSGxQ5uiOgVxe2+BrRkSpjomGyMbTTYQ5eNsAvkGZfosM5
GZQXsHzxPSkt7SIgaO+cetdiy/hVqBec0BM5AX8HIKj1dADAtoYoryN1UucUYXU/chznTGzmfwpO
VRPlQ/L0iV1Op2Vs0tlGeYm7rO7hDC/fRj0IZxU3h1pz4CgCzKO6q7x2FQPE3nlV4ldQFU9V0ZLM
Jt1+P5V1vYfeiSgiCtWQZMwKSGlGUMcMvwDlkJogXVYmKertkb+ziwlbQlI+lbY6gEFKvvNNS7ZM
TBiULfNWPgWbGy0qfv22IcnA4kESSi/kEAEazvXCtMYAFcKJ+y336HgGoT/Q5TeWamr3c1VwALmK
1TzaX5kNuUKY7tDrYo6CO/grRZn+NlEbP40kJqB9tregAcn1Zmsb8RaXVBDmr+zJIkuFxWRifcnt
wVpLUW21Zhh3KowdajH9QS2vNipLdteU52N8iGZW3IBPuY0OqI2wAmKspVbamiqmHym/FNj9oURl
5mOI2IaIfU2Gmm8B3d8icLyNsxihv3zqju3+jNfpACZcoj5FLLMdeL9GQ8YJc+5wcEYJ2VK1O7tu
XfhNTg7pjoY3ee3ladNcsGcO/EJzz8CqsFFWGRwulDvIJEK9kzjGYOck7R3zCVmu2EDxQ2MK8BzD
cO3/yg7dNbxPpex7V4B4libuCrlN5YzARr0UGX1E+ACWIU9YWR0oBpw3kmh86a4QqDEQ/+wgRBuE
75d7d/hdO3t1iCCPtSzkD5REMey4FsDC5KXrcK6AP0EnlPB5wSTNLKanU5MTuLafbYeb83KzLK1X
NRHvETEJM5iUmmwuRZ34qKdB+eoInT1mzrpLU8SMBgqewBksJAxunl/h/C+3f8EnpfOmlUgasHLn
TqmGrjauHcbEElOs5iXkVOum0YHTRj8Ym2ZMinp3/UGC+QnujO0cyCdUnHjKH6En2VoaGQJ5CGyF
2ayxxTH/Uf3SFLxY+5/8Sbin21WLfO3Nw2LmyKsAxxk3heZxoq8DVIXjTiCSqepXX0i4GjDZlDM7
jrOAEqYx1VumV153HN60jKmY5mXRTuuPr5z1mRuMRumdj/5M0jvwoT9qCwjIU6CH4OPRPeMsXPcQ
41b9mZruTk9napwkvtnawxAE041N6AQUe5ny32CC0hFshfpJPiksSsboGhJVnavUJUXHd3QcMAk/
5u6NCdN5Ry2daqmDZiZHJAVMO5+9gWwzhhgElr1k766neojPCogvd2FlevQd/NNBR2v2wIsZQBYc
l7dDQGyMOokEsFtvvlX/X1SdmWniUFveJZ5jc3xe57rOKdLGqAq7dKRZsntGl2q8oVd6wdwaBiV9
GPh3QnkinVkjWKlgtNFJOrqQ4bj2ho9j8YMgOQPfNecAL/GXCaJ0xbdzVghTWCMjsJDgpBPodQiA
HxGxXeXEQDGZQExsgXf4PZNaOe4mH5ej696enrqLEbu/S6ZTHi+6WgJPGmm2DRM9TAybKPoMm/YA
XM65rnp+qpHcQ2vvztYdXaZmp9lPk7tUVjWmEu3CErEGzSuNKt2HNRTX2cQqwcXuNzByHLtUWOIs
HlB+VQbE2/fl01DYTOQhhpGzE7dA5Y/jbVq5ATZO4n9EhxX+oQm4NhSs+FdzGPI3g32sSpnLixmY
r1fQO50dsE/ek6qnSt4qr2vlRMV3XtUoJ5T9s3M+HFEWpEzK7UiDwRmMctr3fpEEmU+rUeGKxCwG
XL5gaZ3oFjGMUB0Xbod3TxSmLJkKQTsK6Ewzwn0LTTF6F+XUL9R4M2ptG5fuIF3YrntOSvIoluTi
8lbW3hdF2hEnqqjvOmtUkm0JoPQeZy9+rilKrXlZfpexv95xN/I56/eN0GU+GLvD0+6YuCR7OyQo
vOwJaxMD0h50JgZKtcKPj8cRm61j/imXbIAp6XfnPQjAwue4LDVfjX+wSjQOpB0FdUMwSFgWZ1N4
MvHBMUHth01IHHnFRN6vYDnne17thGpmoXmq3ts07qNXbQFCdsDL9hNSQ/8rNJFek/v40Dnt1a/T
+XCHbLGxZnRDpG63VogmegTXxQqUh4kPRQIlRCA9coGrkwQ5JZusqAZ8t775lOGin0+QhQ3kQcTU
uEg1tU+Zhe+MGCV9HavQ42v6QA+xCXAs9/TDHtYCR7gYgm4efPN4LKn3IqJdW8mIFKpdV725+x5Q
STusUVJOreutTyRS5oy0LvFOB/2sRnaCNBJif39PbbQmHZyoq8rKYN572ytcFtHwc1SvYwmQxCPd
azJx1iu50N6VmuIkMK7GbE068vCvvyRoEosYYrxh8+3QhyOAkrtgyK3S5gKFMA5bufbJVGlNrjsD
fEtH2QcRGRJnNBZxFh5kcYiPss6fiiQRieM5lHbufrD1Yv6qvWIeBC7iaJd98KoBUh91Hx2L2269
+ax3eYdmBNzEtztO5737LBng5E9NUe4sCdaZxI23u7sZkkq3UDpxrB+Y/uIIOjBBz9D43LFFY+xd
LlWuzP2x/YoRoinnLh+w7lmaAIQ9VKXYrpD80KWUjfQtBpkoqzXXbpqwnKne7EeVUuxikLH6/Tia
To/bDgJCcpiVFVJby8v9UvafQVU57mTt73Q2rlphMwuTCyfBssAOwXEjIYMpxoAQqOqgjqqePKP8
ptDB8NZUYvzjFdseDTAzhLE3NnPLI0H/PTH7/l090Uk2NTNl5AiIgc2euHeMb+KjZeIMj1F8hmkW
WGNrFfMQH4400M8OlefSjL9OJk9AI+9h21htRJTNBsrs+4F+LN3kmTH8zCnABvdn6bl0Qc6Bvaxw
mP369VDADo5W9GnRQD1epfZlxf2I7TXjoxwEioj8uDfmIFqMdE6Le+Y808FpBTEKnmKls13Y9+u8
XZKkaNJz/xGTVm66QBoz/yTXjTLaiU8qX18YzKF3YrTpIw8Mjf3q60DQ4pevi8hTz2xSRQfkDNfk
kz1e0nvDb6jJnJp+KiNlySnB1EI0A0BQ5RbgCUVCqBccPCZVflJObaBfqqA5GCcOjNieyuCfbTcZ
ZAmoZMWsHQejNHuaXEtb/qkLQj5ui9u187MnPtXcQKmHBuOYd/6Oe0FbXh0lDPQZ5axmHV/C9I5F
YPg6BClv8iGI+xC0G3f+nPfDbKoTQw8RVkthUn7N20HiN9G6gRCPQxON+DPSRgzr4tVHJow8po19
lK77M7Y91ZzpEjPOZJvy+6YhD5Tl8RIr6FJT6VEvkgZnm2RI4sXQ6YQ26E7iwH1gzkvQOrLKfsKP
fYKjAxj9u3ycko8yzZ9sZz9zGHNuhU9ZSyytlhFz5Af2Wmtcm5h75B1j8/Zn4BuFAvxBkr3GVLqe
Rx3Nw5uSNvPvMbqeCUssVz/He0I44dCEi9ADu1DHrikTkajXt9SPYRomPVhdn0QZSv9mAT5da3sV
/hNVPpbJBo8HnVnd7yjRQYW/P6T7fVj96L5UDErlPtDSOffA/YUAIEU87QpuMkKGy0gP30hZq3Ou
62UXFeZgGU8u167UlCUOoZ2KnRSK+ka328zwUFEY0oIi0Rba8tY5pU5r5Erte156Fmw7Y+zXe7MO
du2kH51XprKUFibloBVI+ExNF3suDbg5J3wkR9z3zqBnNHLKOz1z+dZnSRfr1iREdn9wBv90ouRb
q7xjC4jUKbf2nFP1A52gsXJyarOzL57oUYwGC6gb16cElsXxdZg9O2YjqM0xWU2OdUvAbCtx+ZtH
hHq2C5HEKcMR2BPu4Z89i3kNspq2+rGp36Cba06nBkLjDJnAQkCaKsRYpuIFMN6RsgelG5Nkd8Ja
DczOxAxGTUO+X/FhQyY9F2nMw5NiM3lWt8NFnozIPpBILr8f6WO0M+behhuZ3reKZqmjT+YDYt9z
VDYZJtHNc1/k/AxHR+BttIVCySHphKmQINWZhbE3sqFq0w9DbEQio3tsskEXUZbi4pcpxH7c8EFy
iGiol7oFlO7dJhaOQ1uLpYqmvDfSNgyrkt6qk20+3Rfqc3HPHuP4dH4FvXf1hYQPlJVlyM1KHmcp
RJyn6RMaAD4hlSHmUbF3JT8V694HR03YrffZ1BuzsUaRN73EZ4bhg8FGq8imH6BVLbRKpN1M7tcZ
dZ0GZv/vjjyzqcm2vDepKpni6brhR9K5xK6ZK/tnJYLlJ3wHOGgsRL/aAjPpyDFjbO11e6ouvyR1
+uxOnnlLlC44XuB/tGZgqBGmR20gYVTw3xpG/vCnNI8F+LkZaLcZzURsfwU0mxSsPiaIjfdih1i4
d12EO+VH3MAVWEHMg6wPKSxTHoEWOUG0ajpbCOt0Eu6yVVWEAXksEcnnnVJ0IbFoBmzD8kC9rTo8
NWX2VT8T2R3ie3C6c+H/ckzAUyk3pB5UVA9O/5eUOocnHZP9hdUYi33dwti0HebuIXYDM47Hk/uU
B+vE8OzxODSEJqYQCwaeSkhu02I6ICYB2igDj2a4CLDPYrJe4WLjo35cVhLM4KprE6FVTaj8UEIg
Yqcz8V1B4JruRrAtuVt1n4EIqIvxjI9ZVbCyx42FR/i6MHXg+2LsS1Z4mUwePwBmetE3N/YiUmku
pzDMGP2UYowc8/XOkmtHA5+r3deGxE0SiQ8vREyS0fIMSnhi7xrscXpXQyvS6DErUrlOrqz5qqru
2WTzOxLGnlslizWjv92sIYQ4UaqY6gZaqk9YQlVuE+jWTQVoXgaJruxPx0hYwNFtBSOWDD57eXLm
DkFGa8ebJN/fSSAe6myOAP4kT+jFyjyCJZ4FAK2EFvkv2kplrmKJReLtuLReDQvQeERqtVINZd7I
74YcWvXsmZTUSqtGFUIuGEWuWIF/OjkaVXeD+AOwr1/MN8hY13Y5vBgChVvR92/JY/RX8/I5dP3u
2T6/+fMJ65l6SdWwZUM3GGNqKKpA+ZaR+2Oy/pB4e0inw6Ybnnp6T7bvz45tNawyZv1F8ZvYZe6f
I5vFGgbetk/PGmvhDD3h0es7369HeFj5FmS2GxlWQNzz4geIwaukpB2fXRPCWNeI9WQowjqWmM+9
lo8KBk2ldMOhgQHvyQpS7IUvnLugk7cAqgEqL+JZDge+jo4JqWGGSujCwwLyCdYOVPOL+QvrFG+y
g/uSPPUFFpvG7uSjB4O9/8WLhmF8OUPvypmM6/jTUEbVyY39aE/G/6aPUkDv3QZXL+YYTxRdqtLW
sNSoZ1nWahJ9EwPtmvEiT+Qzi7qVfPAzuNQjaRHMPREml8ef3uK7TzqMkxIDSJtlcdP6gdTGIjLO
YFHTL0GIPaJKX1X7hborJjMqyrEHHtTcO+i/pl8AQOIMgivPwo0JROdM7rns0WC7AjfDU0gSCBF4
W9Ic8zoPVUcxFFllkkFJS3TVmvIvo+1jnSwRQe9dnOyCsLqqFuuvqFunUzd9bOsjjva23P+yXJ8l
Z/J+kJZz29jSofn95iYXbGzFqM6AF+ftfPIB2N0ClLwrK8NMfk6xltNkdIhcD30YHB8WsTrI9N+c
9HzSrn882/cxHqD+t85vQUAZ0nx3sVZPxZh5cwyQYphajpeAHpB5tjhdVf9k01kb24Ev7e7rKU9w
AYC4QKQBwHd2hEEq21CYjjVMUb5AVfF+rL8wttUcryumWOJJ1yj+yLB2DjRZInV5WMAPXw+6tt71
zeneEnlS53aeyB2FLAsDcpCRmyCv5YEl+aErTjkDe7sBgfMBlMsvCnp5j5BUo6DpJIcfdd/3IMbC
9sEtOkz5ma2RQt/x8Usa2Hkf85bBXa7ruNbvsZilTGiiR/oxTCSGCRJIC9pMb4SUiHaqO30qulJY
c4E9JW3l+7OAEHmxZ5p+sGy4y/c1ZegwjtVi95M8TzEH5l4pxhDEHlIaf+dDdjrI4GuJZFzLsVM/
PrSW6p5+DRClgaUPh6cPj706wt+VqZYnPenRNu71CRhJZkleUFonOa9JfA4njHz70gU7W4hEEi+1
3A5ZKZHVpibQMsrAEUohPcHflnExrDUSkQuBMm9KpeuxbbNn/wWwsDidLQLPRNlv5YmF+PfAFHI8
REjDltmOUr3LTJMTRFQ85s8QyjkgdejdQV6OohI/VTytA3sEGi8vILSoTyTinSGn8lF8bUZMwhbL
jJ+J5eeDMVFvFrcwzloXLsnR3+uT4/iKv9tTyVjo/W/FQ/RVlUpokfgJ0qPZZU2dOOUAi9E8M559
AMaYnA/KhGf0kc/5gyfDL+CwHjhqpZnEPDHatvU4/6hVDkHF6/sWHWZoi0QbFrWX0ye5iLxKyl/c
LETzYIao9ax20IgnOaV4og6AjCGztP3mx1FccWne5ZAcR5sqVqjMmc8NxY2ighuTPOD2y/k4u9xe
BMaIXMHAsUdgogoiSSiWcQDadgQUWoQ0Wrxu5g1CCpMkntPcY4PkI1hkbuiCc1HbFHi7rxmpW/0b
YXnYXPYRXAOHgvMO+wCe91+e2KqU+f/d16RzRMceu1IvHj5jY/QWpAn6AUXRK21GeGSPsczjdeRg
tTE96VoPXL19ZAALCp/5Y+JMnh4+B3Hvk3RQyUsDUZbeFewajlnDpxD4d14y6nQ6oDBzmTXq8CON
QFwNqCaE7HkPVWusi6wMkdnutV1+6+JCPzBy5B8+iqHXTkR+/QelNrD2g0f82eEXGBfKDHDB4Yma
7DvyDWc0yo7bzfHSh/s14Ldt7qt1Cw32ZfYt08JwcE5CLDNRcqZ/q7jPTGJzkH0g2XIViI80UMCB
8SBMYZxtTBpqgITxUuRPT+G40yFCrJxpDjAUP4L8hatO5i3LMDG/Cg7aMfFwxS6HW4O282FvUQ5U
n1f5BaJesQXCFAifcLhiUMWvGf/6FJDK101yPx/9IXQkmBzQTIHUsbTqetIXcx2GDgE+wKh9JTmG
CXJbkgTwPlMnmfct50KZBuEr9RZGKsa0UamAPMWOHxPRBNlsza6JjXNwkrmbD+Cv/jGaJtMjPb/I
416rloPZbm3oP3EoUyXnUIWC4jop+d8qN+4ka4dXIoDSwmQjJfDZmz8eOgJXkYP04IYdbyqBf4xO
JoHiEcmGPmzUgSuIE/hRTh9CiLtHP4Kt/WL8M3Cn0evf7QCglH8ajCq5RcG6sfdiuIoTDSJMxoob
UysIfEFuCQfhvXmR8f27pDGtivYBV+7/F5SvIXojZeTh7JCDUj3y/CMS3HiPWOKkQeiDX35bUZC1
FaX2RL2WnfT5OQ3L9f6AlwJFnINsKdwHAudD1cTceZ9gEa7W7ru1YZ9ZbyWmuJTNQwLCkmnHIJKX
oowVJHHS22UAm7QWHtsXF9qBpxAcBdGNVueddJOaeJ3a1AjfAXBPsfzYz9v5uPxpD7UsR/Cy1GAd
OtW2syCN6J+4VAFN1OHfEnTOFkNBcj/4T1RB+ZUXagdf0hJ5bVtolJOrFTikmqAUtwi8C5S0UDB0
xw8Qh8R1ZiYOvBJv9Z/6EPI3rTp0G7k0NHLFmWckHYiVNIxn8E4Re+zrtkuNbRtpr+1qhHu5vlvE
MELlaxt6berb5GI2k2wDrS7lhKK1kTqqM/GZ+MnyoX7gANLTfgsGZddgiLWZRyfC8C/mTX0NIn/n
7Zxv4n227F9y384FQZznOZuraE0O0pU9SLP+qo/BxdRygnj+GblTQIf0xGmvS7+o+bEPMB5AgiTV
cPcRdy31rHi9AMGnHcR38qIqqcfbq1EFrdHa6Hegb3r27rL0ZPTR07TKk54Gj093M/Ejk2/cD8F0
4Jx3XeDgBh311fU1ASQKbXNPX7jKhTJdHGRlG8RxjbuwxuwJnKoUtYH4ft3b6HY1IDzVLeBSQ7gb
hhVm+ASR+flIwUJ/Lpys6WOfsFoQjxwFW2DmxHyJOJoids/B9dV9NhxNk+qQCZN9uW6bjhlSWI/R
DNTU+ctDqIVG675tGaS5IFrtMpl4CTQdTnMNLg+ViZ5BMpOieGOwJCQIeig+VLW2G/WldIjianeW
dbH2S6ugJNxs8IRP1ipl+mCOd5kpgS2X4MYP/U/FssZzrOyhT++as5tcWio2jY0HkxliOT4iqHbs
6AG4TIcfq43gnVLxbPEBcPdNT72fMDpeBviNDVh1WY34Bs0dGohnibfbGtwA3UH7N+WO4HFPBwyt
GGyYz9pCPqD9DB6S+WgKttgmvY2nNUCtpPcuChfAkAxV9IRBeLM4R302Ip6DL/RvjnrsyGnJt8h7
X8ZsERcdbzOG41GVxUTqtLwbQ3CpnRxRG6FLgDPppQ6sM7DBsoQrqEmipQK1iKWRaO4AoaCUR8FD
dMrPg8rKO0gGHyI2ADid8PIzNz/lSRv8KQj/W0yXiZsJ4zazo1gfAX8vq+/RXsVOYK4aMdGF4/UP
Yw+xG1h966459VroiZy8+JBbmh/vLLp5YTe6S3MPhev3kthwJ7ZXzoPOmbok+dyA4DArFljbjlND
0D4whtAkxgtVbJIbt89fSypSiviWlp0PHcloyM5LgAQaCbRMF2VUIIEqCLQuqvBZVIxyZEjusvso
pBq7oyK/2bnllQQVXrl5kY5v5EVUdQNjTL7+DT14Q80UrqYM87XzcUs9Mgvmc15UeIA4tlieKrmd
4vlTJIRHJNodNbawdTI3beahd71k0ZN2K1ToL8fFCmK+c9ecnV4liQCPkmAtgGTDDKz7+R3LcKNh
YEXlxsulTvS3E3skev4BkgJHLgKx5Vo9vYt5r7zjM/VJeJ/XjUJy3+SpQABxfV1ycOSA9A3OnLUq
D7yNK7XWPecnhk9rDU4mMMmMDhiCXvZ/kfLr922j9ohgThqiUhkaiMf0E6a7vU626/tqpvgTN2Cg
6HG8aYHt4dd50UNFJOdg2mBF6sVzzagTIGBL+qs6suhFnWfcAA9oBFZYRzJj/4aeT4s/bIHB9nm4
S1zEyywK2qVMV/uvkJ0B8s//HWCu3uQUqHUhYaAyWXRyIJdrI8Q2jPAxpwzkyW57wPqtJOBxWZ0U
g1ePYKX+7V5aU5OFPQJKkqgJTQBGoNV7nBe6AjBVaVF0y9Slt9NP5BMVxzoZF5pCOkBeoD6qPB1P
Uw/5AZ8j3M98aZZH4Zsxm9zb7v1OgLtVm4mZlA4cCtXIE/cBABdXtSMBWJD2/KFhusn9qeWNxE4Q
JKpFr89/Ec1k4FRa9TsywLPIQVi0QBwJqjmQEiX00LKX47RX9plh5J5ygaDy0KtCQO6U+edSjLkl
31XkEJorSwKCoObxKMcCOA7JjRrc096lfk2/q+VzswbN5lO+wVFkqgW3Kwv8aqIatzKbFZ3gdKP6
pv3bq/YvOvQtGBJ/IkIyksymKnK83ps1oDueYYVq6HeeE1msfMYeH3NIabzuW/+tpRFdKbNVKawo
vyn7v9TUsE0aFS/phRpx0C81pcbOQ2FQ+86ZB9+fFKLIjSKolilE3AQgmiLbI8i2PFs3vyhpcsPq
HTusHQ2p555XvMzAAmLUYWvDh9KPCnlSjlDt6sPg8WKDu78mm4xeoDGnuCh5u83WjzsYoXSCFHOh
yjj1kVfkhRExRnpneSOeqDPKR1hZAiELQpHRGllrRIK0eRLoy0RbBkCw2FdG6bAsnybYpLKpM6zG
ZFbc49A5+QrTEt8nHgSR4IwINrLOpyM0UvwBHbYTmpn6/yHVLfRB/fAR09OaAdyC6GKrUpQHniyR
j567vs9W8M4QHt0e2hdzFyM9wErdWdEQ/PacpEEXbLWf2mUQok31zMYKQa9P+kgmEqLA5Xu2KlIB
ZDSsSNEBZK2PRLKC6x1SzMZBPeaIjL9G4NWJLPUKEJxZCu+QrMPxlvnwzUswRrRUVqnqXAZUNo36
l+d2pjPJzxs1FgodgAySKhJ8VsThFzvDLuRLQo1Agiw0kM3mDYQ72zz1SXYt0Yb7atwyb4DQ0jWg
bPCX+JZ709Sw1+sOTfye8lnNIroJS5x+Tl8ExxxanIhkq4rKyszWjSMSajYmreMOlE3rSAymQYW5
17C5rJZeo5qAa9uEU1R6Iyijp33Dh+nTTGxH3dmpPE2No638v5zX7SiZcG0MYQcXZXrSOCjfAfjJ
tXnfMdJo1J5p0lVZBHX3iRvwT6B6zQ/1HJy55qy9LB+StiTGM1HqVnOUglSzxQbcyuk+zXJAI8YG
wDUmWKBpfGfcHtmDLr9ueSvkjnIJnun4YwxN6zKRSsBfF5L/9qRdRXU0ZUA4h6IN47yPnknt7ZV7
FnWYKMy9VC6sBJ/YSFDg0HK11cHG7Q0qYPsT1knkPjCmbXYj809/xP2YZhjm0aCNtggmEy2PP8ds
4x4zDsnPgLzRTMu7ooHep7hXKI2snRd12P9b5Hf4m+vbRE9JVLXWewqwu6A+VLi4H21+S2sM49BQ
56JVnoCEb/nJADUbEdJzmwuBNbPPuzo3Qn/kj2dc0NCInGpZiprJ22XXsP67s1zkM151Uo9fOYba
FlsbVJpq++aUfr8AKj6+y+8LqctD0JLiA9bcEm6dl1G7Qb4j5XcjJJ4w9UH2jGz7kbzUr6xNs0Wo
WWzUimSUjaNJIE/eaizcIk6GYMKIGyZzWkVfbUqwzIyBTi424j7BSsi+2JV/qQCPr4lvjZbuFQ7V
wEGb0cikBuvhxh/aEqzdmSEwdjDR1OdExJVfk9rdnh+PUfPUdZdO2qDGZioN2VgPo0/YDIgoUueV
J6aUSl0ECM0VzwcMEe7d9hwr7vVaH4r3KPPfMqB/rCdqCIJRT1SgFVy/UtYvQW4eXLw7gCPCTyGV
mmJ6gIRPDZwEqN2xsYSUyK92Khjd1I6odBuxbgZhW4Flj1hjVUg7O9dOuIXfijfJRU4Bg2L45ibf
Tr1QzlWYu8TZYys3fO2c+2VWMfMugaE5X8iwK0TP6Zuy+B5PWwLsgnahmgw/5e52w4v+WMDe0mu7
3zGZseiIgJzjAnm4lCG3/4murK5L/7/IGl0gtMqg41RZei/ratK+qfkZNoOic4a2iMMDW0rtyigA
dM9Za9hUFALaM0PKuph8/fKVTsgs4MccCt+ApF9S2nJA3EcQIrhRDtZca3Txmu6PNaC/DGHDjG+6
w4I21syNZIDyagEt1gqiuRWc6HAPsLUWFTAaxp39b1bmUtP9+4cx2Sq8tHsNTo78AhdpeqqXPMSr
M7XrrFNPhndu/wVX/+oD9GqJGBFPuldr85P0EX7b3CcaGo38ACMr4G2IeDADM2vczgl1bw4fsGfL
TScKOFMv7CQZ/ohUyiuhVZgxLIBkr5jB/3QFQLyAl0i+6SxOMYfYluGiRVAvZd0suEcTaZB6cnWG
KLUVTrarSyg6bg7Maz6fIbQB2Bzqdm0j9ttXzpzRhPFfDqfLyUAfiaFxklu+71eBQRaKfD/L66d5
iOPBZtce+5WJe37kL0vNAYzJ2500uiLFV5LeGRwo3EY5os288vVly9k7AF1uQgouDuzZ0OePsBOR
uAgYfN+yEEopfcNLyx98znX1xVx8WOOozNDGAU5rhgoC4dY/aDZjjR2/B8y4j3vFz6653qkwkdu7
lP2e1SEJ25V4Z7IIHyaNc4nR++2lFyOb9SqqYkH7Gs+jjShkS99+X4lvBjpsCi5fb2ahuoEEipFn
SDJ81f76R03+8l0AD2zbgmtraVWiHqUt0I4adn+kiXyKP9U6UcNzGRIj+zpRR+MF3r8+63rE1pnr
hiPZe0xgvNmvrhBZpZJxqprH6XG5TbuTtAU8JcIbwJTfXQMwvhRJjnc6j6VkPeGfq9LCVuOM1ShF
ntK7bpbfeBQN9qpkeHHn88NZ0k0eehU5fFYdztoi7WtBW6y7whJqHJNQXOrxYlicrluNwXVv16DI
DpbZdOfoDOQrrzFXvFyW9pVHQa4c7bAIVliHurYWkdqIW4NRnzHfWJ/PvlL6yXqGREg1us6FGOmd
S5O1JyAul9CCFDGbdRSD5WLCa8SVi6zNjHIbL7ri+AqmuT4yZJd1efDq+9ACr5x3e8fMMxoUKMzs
8lzLh1lhz9OOJhYbfMBnCPHcsOrj0nT3II8xwqopl5ol2orgE0sBWG9rSih+BtVURtoOmE/gkuxk
1v3aIb1j0zP4UMY6G87wNe1nGeAlhK8c1V89rSpIi37ui7jd3wGECVA1rU8UI5N2/7ulVOWQKJvC
ojOFwJsT9aKPPAHlbN9DrI3QQgTIl4UviPX78uULNfI12dyUhP8hXp3CdZVRB6kBnETh1zZZHu9b
8TdlLmfHyPxSN4ndOMczPUpUIvUqKqK1FmfFNcIQsAnfdtRRbadBn53gnyrXGxpigckOQy3gEral
zbxWmgjwdkB/HAQ6K7/fgNnn/BwgaSeJmHO9SJMk0rSbnyfsRtLktbbJ8tRr9NaVhM1fq72ThCCR
KKHszMr2EER0N3f4WCqpFvMZmVXLdVPxmgcI2nHu/Iafuz5isAE4s23SgiHwZDk6Ag8wNz490s1h
B2N1lj3LWlrJdrTmVhA2WQaPpM6pTCHsSCsE7XOJXaaMvkChdW0LD4XpsATgpEqyHA07xXVp10+W
ZECASnoOuk5674rGyTkXojd0MpwxYk/MD1dr5MN9Oxa/NBtj7ErFxjWnIETxX20qbgkIlkpn0Gp9
JZH3Ar+cKKMm4E52D6kvQULD+SmWm3evusEOYHzomMWrKVwpH3LWKvq1ixngwnIQI7HodAiOidep
WbqwqYuiIaKS/nNsmZTxU0xXk8JibHWS3hpRel38AFWLt+PTZWDMC5T9kbwpm2ICT0hm0tagmQNE
68MYe+DVOg0UEsr5iajNnX4Aj4AeQRW0yg1HCT3noEmB7SlyxZKXjfIMOQRzwmrcORBAimeylsak
kSceBRlER4MxqNpBGY60lUWcTZJZEQ+ZDzF1TgDJmr9u+1XBVYZHMMe2ErQk2Q0FYH3430zwALrd
qL5T7p1QbWaalrmjsYDkUuQVI5YvcVxmAOPzrUrkgIhyQXDKW7MXqpvLaYYSpGDfbQtSvowaYzYO
OiT8TF40asuq/Wj7h5YTrce4No2uHEuGLnbm3I9QC6tviCm9O1XPMO7Xfs5QbXDY2+2xszXvCsis
DyDvCI/5r4d6onboEBpT594Ht7ZsXYbh8Jg39RRtpmGc4qdo8Rjt4bGX1QDjOmk4ZzRX5yMsSzm4
4UGhHP37m3Sxla4+kJyY7fNd+ywY6OUw43OKRkVWhlSv/nTEsu3mo8Qr4RaTai5bqVU83Dxpn0XX
6OXHKBP/DA0r6m3+A7b2pf6127jk9qXvEOADZkBaINhpKvZamCowAt6jCmzdH7QL02JG8Zloaszn
solmbuFwT/olpGOrgfReAsa4w6Oc/JTXisFM2HMv1hZyR9jLXFMYcuUWnmP+efD8fDHkr4XlM7Xg
CshtsMpWygwRdWbh15e/rIJ/4vylsZ9vtCLm7J8TO/F7/9KNUQPbzr6Gioqc9YLS6k9dG+1Xt/Z7
X/7SX6Cw8lQzv3pNGShaBJljBZexiDJ2eG933JNHjd6FnI5Jb0VxQrFepQgFymJ4HdGO8Lf+hkxW
z6l+59uhGj1bUj5mj+mVlddqZdq26zfYlK8wKssZBt1Djgo2YWyntKvtRLl95dO82hUYu4QYZyIQ
lgTyCLhTLG+dblJcAbMkTQMymhI3DW7LuxAF8cCe29tp5vVZLo/N9CE4oZk+x8QBYHoXCWTOCuD4
FyCCXM/ejKX2Fy2oNOgUDMGpdFjU7Ij7zU1mPWkgTCHYi2nsAb6JP8sdD7kWLXmU3fvYy7UEWHXv
A2Zy0EQ5wMp30+ENeTnmHB25iTns7KY8LfvLhs8ZwtlTVSIImLHXIkFo2l3TvumtWDaKucyJU4if
TlMyfFyhjKpioC9SxiNt6wpEbPHfbHdLWTj70PkxdlAPX8S96vyUIAJ/4PSFWSuOq6oKdD3GFfht
+iScWvMRWFOkwBo1YyC6f9n775qrtsyeDCVfWDfPWX+sX2wLszjm2LMKSwPWzKaeLuYqqOLn5GJI
1oaXqjhywIEsRm2azJY1nPE9F9YUcVf+Yj4HjUGeTxKp38FFTTkYWElJpjA1abbClIUy1VPaf8XA
wfTINOeRvVMtiDl3rgpclrEk4oBKInsKqrOKCOZsTAsSlKlHvi92aOYqOKNUrEN1BzBoCsdDHqaa
rFx2Unj+Yll/oeNgV0yTRSiGpDHcHu0WDeaGVIYZdBEWIEsMmmTb13msbfQV+0HG8TfxE+0MAzZU
miBOdIxo0aBtVXWmHftBP6nl2upCOvicPinB2/NLlEsns0e8lWKvF/2RXdnHXimrN+xfX5HB2K3N
RbGVDCXuHJpFlVh5JAe//JFBNkRneBweHb2JzNy2zQo1SHaNUYXvJE/tMxdPBbs6VZTeoXTW/Int
EufM2HfcL6Cx2d/tfhWTJ5Kv1dZetpp/7tdRNbdLn/hmCUdJfOlVkvQzWGOUDqXorwXAm8vzvDNr
BPh9S7yM1Cldb/9Y0Qk0zRrgY8GbgDZtc8FTliqXBOCW+E3th+UiwliEy5+kE8Drv8hQWZnbIazN
EDDkEmlPqKNSh3KqOoXEVwqr9mkWvdEB5NNg6aBcYkgFGcsPThHCBr0ltrWjTMhEyShit9n9eGUy
zZVOlmOK3FkZQIrBsIX4Fw7sY5oaWcTafkEnKwtsExfo6d9Zzx5Qqz58fSMSbvxiW8Uy0V8XE0Bl
iRqL5aTKSPsIJJ6Jxb6z9TmmJK3XjwGj8SSqUt49b/DT+CL5LianRtcSsfnkMtgzBjNYDJvLQK7W
/N5MJ+CE2U5yosJxdq/SROfkOWj6AsVHtXZjwWUZG16AguT+t3Ob+7kNH85JTg75/X5K5kddSwY8
0DgbgYxRxH/vn3Zs61CPcwCsQdIcLnEuv6lwKxlJKt1YugwMBYUG03V9FFh7lTJi9ZKW6e3ZzDK0
iyZ+gxIORJpq7xNijx2n8GPaagieIucRA8E29YP8jPyERo8nhrUBWB7dhTug0+9xL7rnT7ZK9gow
nq9HSgfhfhueWoC2JMhM7kHHZwcyRXf6ZsAFXYQ3YFyZ4X9R16YQUl3tLz0PvrRmoe1tvW0lS+5i
duAoWSwNTXAEE7lz0VJ4QKdgfP/MtS1FyxvKZYtAmYUsoSCXwggGH/+gPIhaDnRrOvgHN/9qKBpx
enLoVUiQxAwdFt0jS2GoqbTDdg+9WCNSBKHVZHmwNQYaRpHn6LyCAYaDiq0/k7nxlYH6yJVafntc
ZaqGdFmrAOuNUVVN74oaKEgUSR1Z+HIhvUbKmh3vyqSAoj4dZQWsFwQtqxCypuSHQRolCP+km4H/
pDe8IZ7gcFPXCp2OOucJdq1qbCHVuwXrZeAwMAJEfkUM0BlSMzeJl5nrgj45SfYayuN8Lwd69blG
8Mz9AZza+oxxfnmR3igTyp2BweIbIYoYRXTO9/BHV2GS1O/FQ2x9nIWCEZY0loj+R3hbluGtpbxF
qGEP9dJdPxYqixlsHiIBgitIgxr8/9V97tKHQNmxBu1PVmPLXBDSedsTdMneJcyhB71ShFf98HV0
LCDuc2MjuIi7W4K0zIpez0Q7YVhHMxd7EKzYbYvkOYZZ4CR3Ct3KMuxRSkpxLLOomjyuOK5sbu+F
5cwlS6EbsU/X4fr+sY3xfQW5ZEbRGXUO8UxUYXFlX3zDsx9FQzK/OnFpZriws91A7a17V3kxq7Y5
albD2da4SWRGHjh//GalxnO88WWlJZ0fKcySa09FRRj6oiOLq2HMWeCCS4jw1jVA+H7ndfJRLO7I
/hkraLgOfrEbapmImx9QDxnk/IyRkG0dw2W/W+gJuK4+sl+TRAbwX4hRmutYTaa0GUF6xM5lTgHn
EAve+GgI2QyD+IHKGIfevERuPhdG76h+wJu45gEId+NKJ5DbTmnPo4lSzTbJvrDcoadhdy61h5F3
70SvuFAPSbi0MGsjybGiAq3/QkHdiIY4KiU2EYP4H7Z4GAuaoP7CdU7M82qec9fiONehgL7UtnKD
9w2hUhFC97XIQ8HwNtMF0RkU2/E7ln5g+vDeTli05A9o4zMjXPe5/Sr8Mp2m01/y0pSyHUrFki0s
AL8JtBh2ydYuQqBOwVYWuXAiZmxQ5SjL8KXxCWdkxFZOMLDnEUBuoWXf5wNly6Se1c8bXbwNX1EE
WkyhSThICrY+aGWWiAtPjo2QIybQGFaF9vmxqIthfF01u0uaFtU+PHZvueKiHKlSwM8v7onmFqP7
m6mTX9kXYxBJBRCxoLHXE8wWkPQg468inz6s7vFQ9wEf16VO6ufSowmwC8Vbo2ZLbAJr0+10Cf8+
Au6KFqjR5fNTEkotrJkJAvWh+i1ih8Djr/EiOOYX1x/dib7RT71mLcyuKmdrni3w1yjaXWgOsfQO
dhanbHb/8nVGlBfkxVrXnVPzGSD1uSu8Ln1pXjGsFOFnUy33MJybLrpIutGaWfHqGAfsFovPo5R8
zRboBs9QXkpnB3kSotJz3QUVObrSXWYWfCvTQYygEshwRcApTaa70BqVI6xN4YzYepkVyaWf2S/l
7c2wV71rhPJCtyu2GdeaWxcZWWLRqL1DUgEk9iSsJh9EJgCHrn/qMck735rtEhNaQYuULvhWGNPk
RA1lOSWuxndm9tDdOgG47GX+2YHRJNBuCMOAWWLBt0yvXdoCmA/6IjS0IZ2Zr7RaUZhFSvJY0BLM
nqs1pAV5rWAxf240uywzU9WIDcrY33VC3CLwQL/v3wGQlHwf8mCxiEmMSPVW/TF0RVm6x1LxGCv6
CLKf9fIZsoOQ6n8V3MwhvStC/+5IRMPubbaci580jQkjncZjZvQMej3+hGIcxGZNab28gK/me6Si
F/pcpHJ5vTxJLhmhTwCg4OjcQ8yQhAJwV6o4YE7uratJgfbBrfVd0SH2NU/2D7G9tVcJTLTmVu/X
o3T4xfXFcTSg8yBGc5ODm5HzwN+SFEr8Wt0O78qhEwoIbFhrt4mga7N8c4yuBQw5uxZJpTkhEzr/
w9RWNve2r1UC8H2ajxK0wpHj5OYEDvBOJnkWUKhuqwyylYy5AShyzv+qyIb+JYRc1x69wTCUtRl4
gUYhdD78FdPXM2X07InwYKZ5UBiVsyHfCThIB8VCdv78gAKsuTWzW69UKdSx+FHlv08LAvEwfkl9
j5P6DbRSerXSUkiy1wN94WsjxS4EE1B4ckVzdaSXewMuINvoromW1wUdszW+qo+W74VZ+83dK03I
ykHpPgVOwcWzGPontcMhmQnIcgp0jIgDlIGUjEpyt+4n1lpwIyrRUo+5luIEd/Ax3oBb3CGP1CFS
gOtdVWFs9ZDLFNSQL99sP79QFcioYhZg1fBmXf7x0fDda1I3wFuwdAimF1axT9hHjGv9LYqj810P
/bToiIVWyGTqTtScwPSdwBUsir896s6C3nbc33GqVOcF2LFphcDXkTR/M5RqcUoz1T0XX8hEHkho
jr7M0ILv+pAbKFneBowxZY4+S1Od6E9TMQIlPWJPr+9Mg3UyIiXePqvSA6Lgf45e+4ztLfybJxpV
MDiYKL2PN5HmBlS61fpnjZkXbjoMOmzlzzdrysMYJHGpyhBUxUuoFYMaySm4uEcAWhSquT7tKNng
ggeMxAA++jCIOw59+DFsv+PUf9Y/xV6EWhDrFTfd9Cl+lGPZT+mhVnYlAk18hVR/juctoYf/qcO5
U1oa7y0x80OFKFuEqwFNRyLVuXcgN4BaMaucXXLsikhNAcDczYNicQxPo8iI0UUsdn4lGknBIJpP
Rk7ESH4jdym7Nbci3RWSwhKIe2/pB1x4LKguu4M7u56XLtC8WzpJAuWcAjySUztpE906KT1YJwq+
k7Il3nNHtUFzHvozWBb7gUHtCPuQoFDla0htTbuqvr7/mHeTSBL/u168HdJLe68y0s1xgt3nTAqK
+d9FYKhIcx20B19FcAP10ok9DhV0FE4fb6tmbbtcglueRccAbDR/+G0kPvMMHEv+ujqJQ487nAp7
jxqCIv3COpELG5dBaQwtQt/j0+s66WIt1fPGSdfGZUWGnuWbxBdR1L8gAkhjxlR502Qh1OObJdn6
1BoL2KNTQY18Gnfp9ZltikMojJVI6Xbes6W7rc4JPXY0CKsCDWDrhDFcgKdnIGOtp7Pi+1ZNZ+Qd
eRq+UbJDqWLq9dsxB/FR8V8gDZ8nb/eOL4xNOUKLjYApQRcKe/6k/LVvq2AcRs59e4tRky8WD6Ze
OIFh7eEC9yyxe7FRhCVRpIQbvP4p6Tkmx3u5BjpfqvRKgq7sx19uzyHzZgNpa+pFB1sQD/tcRq6v
WFYiIthQ3hseMw6wFdHXAp8+S8J4dj27WSIhH9tILUQgL8i24d3mgo3WZwS5dNh34W0/aF2a4ZY7
r7798vQlwhSq87CWFnDJu9TEyCOIzlmZjjCTZjWtKRpX9LiQRO+0N6mt7HhK7ICvOyABlBRumBx6
uY5CMWXMB+mxvtAa948er8uoSXQyifg2pqV1jSwOza40q6hLKwOGzJGFY3EahULzacaBozFll6r9
BlFbHas3zp8347/VRz9Ef/MBPjzBRkZ2zhrZjzcAVLE/ths/iK9CHH9BN+ck+dgUZouEIUsFQp+j
C2QLIAjRRU/jY/I7DfB5qe5e93oYPdcl7bbqdhp23TGYJ+nCD+3Q+Qge7ROCAcPsVExwZZEVu6ho
EGBHTC/K858deMCXORW2f1DbFY5lawlIff4RCuF9pY8sUgkqun00jQSaNH8TQV9BleWRcEqLuezo
BEC0V0jvXQgLa6PAEhHraaLXiuuy6da/aZNnXs3TSKvQ8WafgasQ488F7lYMjE7ZpLWsxQTYiESI
7MLvPo1EfvWmj62vOth0+uMwbWEBvYh0QogMadjhWMVuCYVCiFqhM6LlFhSvsbLzgcWhvXY2Ox5u
Ta3y8jMqsRUpEPs7YOdOEDYS6bN6fFMOyTzSqftDs3nn5a1fX24KFcYLwxADeL7eO6tUDrg4YMj6
YXnRGm4Z3TJIj3B8ILq/CBj0oJezxAo+mtqjBIBDQU3zG9Pq1ktjQTPHME410cUQAGbVB/lvEo+F
sRYK2Uc5Btx6WzSVVI1i7sWuG1HzZAr8hTzt8Bd+pUGWJkHf1KeiIikwqhU82q7sKhFT5C2hsBRK
SNUJy09F+2ecl0DrP5f1rI+lzP7PO7ArjH9YltmH3GAXPsBsdO11GVs+emSb69l1JWWygzxuMiRM
SLgNREY+4LtqHCE2GwqN7hELI4HRNrKZ8h9wE5M28NBa4IOLBNgKjYjgJIOZy7t4YzZvr6RGMJrl
Un3vPqm6AcLt0qyTFB+ZUXrxEpV/NGrTVqq1d1KDCS/CWG5igIkMQncE3/lxyax9TMd8pHMzhefW
u/OALbdfGDKnrncSBueWmgTS/b5P6GxAHj/NfLWqnSI1O7+lQCzoLBi20NG9nx5JDYhmzFETHi2w
+H9SsJhQLcsL/Hof+8DTduVlWcRFjGIrJjHDZQkujpEouCaqWQvnY6yEUZZk3DYDJHZw5AWQoBHE
tEVtTNCC8TadKhWSsH4EMG7LtZKjS1ywQY5Ak8fFrmLYx0eDMvviwoFhsKWp+kslyyW/I404Dhbr
rLWCf9PpbDKTqFeG4gByN6/sgipTIP89oWQwIvsofHI+H4I46sFCsDCM2u+UAI0Bl0+f841O4/r5
yy9NUXnofnGd9QxPzRjq9XL9HN+qiHlXRU86KhHDVAFCcWfdmxSNkyUtRVtxMXPHXdlSEKDCQvAZ
3JnB6bJnplH+hjJfuPV6to15eTNFIpIbAk4l5xq6wfOXszyw5VtuM+LNemexCM8jamU01wRzvhlR
h2sFGQ4xBxx32+m9z2UGSE/LEQLlQzwAwZ9bZlSvgQ9/7xdA5mr+UoQZwWB/hoASSDlbLJliO323
EUW8jWtAZTR1hvAg/6fmWJ2pFAgpKZK3GF8xMIHau+QDE6cEz8dEnv1d5U2kOina5iaHJ3LcfpBC
77paYUgj7EqPa3u+HY59Syj177TC2sugVAG7PwBnX8vWczgjBDJCifD01I6nW6Wi7+NGFbhZ+qL2
dcyuRZ6fOAAaFP92wuSrObPyxa7h2AtjboOy9kiA/n3hRYvRUwgL2vmh/sC0xJwrZCgNYubU6WQJ
ek2u1oyymgMF31Ey+H/cnlidNRhDozCUgAYvHhaG4pYAHJvJos7RFO4Wxcu+v2WKWzFTtp3I8RTx
IvucpPTtQHk+VP+mq51QZoWs2CP5BvvQskRxU8ShJC/uOWJOdDlN+RGrWArV4O/4IwNERRT4ZR4l
09wUv+QY/8uGBO0UzkPrNT7YGyc9JzE9Mad8F4hoydIaggi14i6DOgW+4Ulie8jTLWed1dveo+MF
8sUnuoPa/Sy2lUeEyzsNYnmZyuNS+TG8yOhEj9UUK6lxHnLaaG+VvH2ZXcoMYI4OEpAIQuPNV7YA
2snqNjUADCMVfpBoHRUavwnUPFCdnbYY3o5jMtY4fQEHPNR11uK6drBLQJH3V1Law76YjD8CzNvt
Ew85mDWPRZP8ckCGHNvz6j6YYUmu1tnfB1rU8X00G/7VQ970C299F5Gg9itT2GXeFomoR5k0NQ+h
U3nHVSIaxHJeB0Eb7C8WG5fytJVrl5ust2osWb60Ru60OiTlUu5AvoW9BXOlR7fgHQcWUXFxFZME
1vygKZsaRn0KOtyX2uLJkcAwwy0Bqwms7XV3g1dhTM2tOt4nQmy9Vt+9v9VRPkwaANLp8zE66Lve
yRa0VyFkzEYlvbtXNt2fcJwDyGm0lZl6w8gZYrONPjbrxK5qSjqDgP4+UwrT0GTwbLO7CpiOL9L0
akjtgMDiRl/Gn0C0wr8/iTKk1FJnWE6qGqG0CvwKbU1S4PEu+j3qQtHGQt/KteOb89aVp0SxOpJL
wQRCh1QXIZB49s3ZEnLCh1U0A0LIDgCVL8qlgXGEJZcuEnNwc4cTSw7WUayVODwVCe569hGMhGS4
PRIO8aPzv0h76R4ZLkc7m4C29ghyp3C2PqWwOY4jTM6+bvtbmUEzEm25ESG59Joaq/9MWAvU3h6x
ks92EF8sMawBGP1d+AFpZsN73K8+qYjn5HIKdIzyf+X2ZNyAgXrzq0XMbp5Sd8f7i22Vu5iLO59/
NPNirGyPIBkyG8uH/IbhTqm8w+P3VghM0CmqMdJV6+n6RxCrKgiIw0hdYBhXj1Kf/Fki00ss1eBG
Awvv8kAFz4LNICnMOCb/3zIZNx7Ha/etFs+rOJxHsXdmrTqljeSz+O0PTI0nxh9fyA+Kctox1kNL
tJz07r4apFLEVSTdp7DGGoo075yVZihnnoDKm4WijCEOhXFOt8BFtWbKyOPOAnb498oaVpqtFlZJ
+OjULf28IBnvNoQRJoLifMDdHodD33zedOnTZZUAWJ1vuMAdAOJvobgyxJCLJBlPimjRcY8C0+Sg
iLD0YRqvXeV8e43AqBejwIbChuudl3EbaAzua32OqLJx1l6ctmt0/XqT7XBy4ZJVFH2mcrWP0kQC
SiFJDEs1gJHkhb3pl9eAMkc2fSNcrSR8XlbJvJ0Tb3b/XdcNU/v3D5PiNMi6NvdfNk7/n1df/d2F
7ALpyCX7zmJ60Fe6KZPsIgrba36QDl8tLkuYRh8DjnV5kb9HnkzckvSLLzgYCu0MDS9kNeLBXqbK
ZEb8L42v+OQBTJTrMV3Ds6s0H/qIEImGHwSUYGyTSI1CIPYCOYP/1zjlpZNgk0s82yRPr8tovHwC
gGz2cpWgsAs9E2hcijL/M4gl6uHpclUoTR8OK2K1YVMgqnbsi6U6m+0aZc0o/4v2jRxIs3f3B4BZ
KsWCFH4x6Ct1IW/nNkrSOutISSLNxTUWzbVwfJXrBdQjLm+/HUBJfY0C94o38WOvAqS4oZ0Nv8V7
wdiUfMv0D2ke+GG6MKDO7k6zJv8srL12fYBVDzFupbwqv9DcarsNDki91YtZC4ff2tusYsGz4pk9
N5DPCkw3FoCV63pIwyTp0n6XfrO1ixxksWqC4yoq4ineKi5L834J1XsonpKDW8rh01LeLtfobflH
yDB6qGAksBbxDW000aaRIuJ0wQmfzZzHebL7Szu0UZIP4R2GJP7uSA5a3h9XoKT3AWdaSX/oTjMA
W3CmdxjG37sKK3YgmAdbdetlg1yWQBwnzXGOS5UshtILs7oE3DXgUir1FUeQDEw+NHAy5U3PQGtt
GIPrZIfMeCiZOivG1UjZ3bQ4+HyfESqu0D6JK2cPbjr0ByAdZKbF4uVxgtmXdPqmu5ZoLAKPLLda
aLGiAqWpmTskqu10dCSKBdOWIoners81fghdOb4T6bl9cWi2e0zFxSaskQ4LHEqd8/vTftWDFd+J
tDiOW1pe1XugabfxMCGQLdIf2ptYIeyP6S9ess01h1JH5K8AGErZpCb1rXP3CjHh4EoIp5AjZcqV
e8vWA+T9d07FP9/tXR/M4MN8SYbEdPl8/mBcmm+gcf31pTol9AqgaEBc/PFi3t8i4CBUbccWrDeu
lMder7NKaSnzIv7j03QXUFo0uX4Seux/pBK7+/WqFjStmJ60YxTPaFL7wLH2DryMBDLq4xSZ0dux
aJpvNoWmjm1oi+NQmpGbkIhGsYxuOEDH+LXAUvUNAFhOAhqIevPkCtE+bwlb8m/DXdVgtrqXGF5m
pgf4lJC2A+6dxrC44yrDWFht8bszPBKBNU+P5cPvZRaK9G17CEL3OThVtWPjJ6kZyZfMGs4DIDp0
SoUaNaZv4ozJq5p38vd4QU8mecbxalSlQYp2BYZ9TiPDemEH8EjvCel3JuJoLNSJCukFrFA0yl9x
BaDfn1EZnFehXQiSVvg32IEM2dGkTpbztk/Z9GyvHv0hRqcYvaf6D7wjvgE2b9ej10ZSUmcn/ial
Tqzrdkcph3mvFMzq6f79J42hfMs/1JkF43gZrJ6cxRMr5u/QSH7Bj3CJ1cmcVP0TkLsnZHgCXR2O
ZuBYDd4v4CvqHKyHdZi4uWoWrj1Tt+XIdqzmPWdhADRk/9dcoDLCQ2Fr2dJtVszMwuWlY3XS4krP
kqrnukJ5VP/3ZJrXEW6uKLMiso0qi9iyCghGcmv6fTD2HvXWw675bt/uLfeUlGSe9/whhj4NOqje
dnKQyGtfAxkYPaFRIVJwzdphbJPCBVYUgHbGO4M9Qw0QPaEq33+MZ6L57F9VNdRbV3GhfhhwoQg6
xGf49BzloxUMd4wg9/plmZPDbHD4qbCYEIEGIPk+fdxZ+jGZyHMgu1IuQ8Peh5wqqf9Wx22h3e34
6amFS5HUEmXmVPDEyxtUR7xiGLqqRPs4FD+91h8GxjUljNGHdCVAC2riwTOXWj+wa5dp0YrcLhCV
lHdPbRibtCnTAnJzXLv3ClCb5urt+YvYgyB+34zT7R8639d3/8fZJRTKzgSspxcO2yTEU5ZQClZH
xBrOLZF6iBDmwQF/i5K3BFKZ860x6LS8iCcyiWSQ8UZgIYu29il0PVPIM3tfcYClSS5Tguy7uzpY
+wxMKbjK+cEjvJNTm/bvUJwRK9KxcMdXmJgnTv8UdaU9slMEHBP4GhiLRG19O6cpsPeQpT07pCDX
y156V+xFNBcxXFWNnkK2meQRj8+XvdKz3EfZWyOruOpMU/m6wiQouUBSAbjX/5O56pmpwpYHDNgb
WpFef3uqCNTXIRsrG0MeYRMqC46CA1YNKkhlF7nXigY7ilzR3i7M6ih95dngt8Z/nXWjDVxRTYZT
GbE1EadUmpi+iqPbMyz12la2khooctKtrXXvJ7zzOSs1X8n6hiamuJa9YKArvllXV6/ZbskDcq4W
QwxB8ysK7uNInnM9TaNMMPThtTBy6IgQjqs6d4a6LnEfAIMbTwqEGcQy3vOhr2VOXMoOKO6Q+RVo
a2QlcBerLqTLUpp/hCBsCrKu+hcMmlc8LPcs0YIivHgYY6zk9lDKARWQUdARKiHHKqWl2yQLnqiH
nIomQ/WO+ygTcZEVohDkkU2bbd+QLycUtEr+o8yrZwvrYLST8eSZa3TSLRBXD/FvCAj3RI1jcD0r
sKSA+UP0X5oh0cvNQxaOyoUyNaBbJ1x1Hpjs83Gwt3UGxtN0fv6Ih1OTONqbpm4M7AsfPSTvGDfw
66d9dC6MAqUJVaU5wiwu8gd0m09JKQzYYadZ0uc8C5+gKrec4w6aC7dGqvSWJiSpk7fZ/aZ/XFI1
7piNCj2TYfbTqL+ltan3zZaTaXVCPockcnagn9rI9RTqvF5Od67ixL5xKUB9NJQZooSq6sxReYPK
t9s7N/8vfUzLxbno1YoCRpI+52TembnpeVAkgMOQ9eaVwGvGHYH0OsgrhO4Rowxb9jXyzuhgUNMe
bjOuYXyYzVREfFEi38pg7lAKhIXgeDmQbMeAiw529dJv+alRqFAfKuqCsWqm9kYwa2twjlih2p/m
pWqqaFZ/biGyihnAl4BrkBwj1X1vzzn5IodXX5w1x/sKDCnzBri/lR+dNOTOXGF03G2DeEMNZnYt
n70IEwYlNIDW2Cfc4b0+/bnYe045nG3f2PniS6dX2M+clM47+gW2kmqzcpmwHIEotklQfYRW/kMR
yEjNrWs7YS3th4eLsuFG4FSS2xdw4rXnapgvPJMMtW0HhEOFF1pTEFYFVCSKYz/QvExi4yL0LkJX
aoGpy7CuMUChn/4zU0zuLiD2MAmKd8Rd2vNeMpCpFsai/kNA8GBe2MqDxk3s6JuuZuGb5n082rI2
cacRn2jQPyPsXY5tawF2NvS7K2u6zLYH6vJ9XUUPefWZpg1tptDtMv7awGtzcgDzjGJ0HeGPFxWb
+OuhwVwsKc1eHEsjS6U3CbTjBWrJt530HUbD5FJG/+MSvdHG1bR9upb8Rs+R2Tw4rGzRz12m9ECM
Ih+7i2+PB4H5R1HvcfUSGQBs8Y20LKNy2fnOBDtgIbmvgUuaxGcpELnfB70w8Hr4A3xCr/4DbbGv
b0PR/ZOuuK9hQoqxXjTNO0kfYdTG+0zpqguchSiGDhmSf2dWt05UvJdijxWNHlW4lwWDcdFFkadB
9qfS/7/UiyyX2a4ew1kvIwn13auchStP6BlF1eOpn/nYDuluk/ZVyF8Hq4WpznTjoblFtwS/xsAh
PUDwfwgVXZOnyo9+zheO6yhrEF2AeqhIr+7jBjiRJnwf5db5Zg12wpFC2oKuBT1ynLpcvybRf7/9
meNyOFPrEkvVa0AuK81/7bg7x+xQNZemoq05hWQ2AQHYY8AGxuobkIkg9HPvdC0TK98ImWOKUgXr
pFaSQFH/JyavA2w/7IKR/ovIbWV4lr6iWQyuND9lyf8E3nUerdrCq9R7DDHiJoRbWsTk5b1aXeEF
YKsKaXTiLJPvsEjkAVUWHTcPpZIp8EIPROugckAs3t2PHcX0QkvNytq9AcZN9zvcOCxgd8wHhQhy
2TL8wts4wqhWJ5D3GtVQ7dfex4QtSWYoETgv30TrqC+n7+yNfGJBiJqK2xnA7LIggTGwc7vsOBdJ
Rg/XlKqtWbL6Pn4Sqy1NuFNinCDTaos2PUW018feGga9+gIIaFFT8igRQ5wIonmAej9av+0ioeki
n7On9ruxjE8XySAb0T7+NjJaDCFcPwLI0UNzXaibl/faHJjS/j8BqWKWATxQcCtyzBhff8hTb5WB
KBktggGTjQSo6VW7/GYgCk+eZLYaDydDf98TARLX4B8vlcuj5D1nmhcHhEAnoY5jAKoG8yTkWadD
rskXusEapEj8gSE19C23QHYEjnVTTr36RbMyFC6BjtfFDuc4LkNrNEMS+KyVjAN2mpmCZSMCymRQ
BzJkkZyJ32JXcLgEAfO8j5nT/FErgvxr3FDY+m/qhEN5fTqPcqH1D0vIc1kTyqUos2vPNst5AOEj
cjOKsxMFMTfJyr5a+/d3cyWfX2jsoIKCJzd+2Azt9AlEGEusjXT3tPIhJD8pfuDlkjjAXnM1ZDgG
u3toBnOMFGbKdy+iNJmjtlRkM2rIdzi64KXbIHXDcd/X8O8GB0loHPPewvyWdXAA5PxBM1bi4QgI
zsHa9P2u5F46vNeq0SeVvlBZBM56T0WhqyTkU4kZs51uiE4m/tIgJaergT5upSW5P1GJvTx0wFjv
7W1juklpNy7zmV+jmfrTIePSjfwFzSIvBAI0vSFEkY855h+nwYM7uY32XBAGMb8je/t916rTiZx2
CR/ZKd3Q1F06qBre2cZgYPthWjZuM2fUrX2fpLTkA0sG4ePoEZWOBW+8HrZn2KnSxc9+t8j3f8Hc
DaDkYAaYLh73/ctuAH8dUhWOkVuThKBqFO1JkyqTUJxLWsbopqlSQaHFMe61Qd098koJ1U36rXu5
Qw9DgIR1ItDWibgNajZGIOd+AxZdjPzoqaMpURjGMk+cwLQ8+2MiFhPgADOk9GdXPS/zScyJc9Iq
1AQFHwQ6eMhx3omNMKNrjj/VKlYwElEfjHl4P+1qpjvYRUOH8+ZDYuZXpJ0tJSv0wuNBU5jOuhUl
nbtOQqh6Zrfb5UYZmDOZOJxhharKSsygNlxTLD72529YuOXd3emWB8+i4nvs+R8jfR+CUu2O6qH+
rUMUT6c2+r7o3HGRghkG7D0iA4j/Qy+MjLpxwTxmjsz1NyQBmDfquUuRMrgYZPa89S7vb5loFx1i
ze3e5DoSrowIoz2i7iR339NANBFdI5xsafDru+2ntTJwN8fU+Y32RHzD671PhBPQyC5JGQCxj8+N
QgP6iJNCzkAsIExh7fV3h4b/TgXkWlG7bspeL8RSugh7nHkRvpbiLTN38ard3+Xn8nRr6FYEAMnU
uTvF9cNmgAh7aXCHYS+KrctxIs3DjunMbHofroMbwRhyA5nI/hbpcwtILMsOHrF8wwVTNK5fjIcf
zfpUS+PkQPH7JXGF6ZeHmZpK1Ea4bUQnqfgyazCQo7iDs4zOjABwQSQJ6gFpgKHgGZOFNkgMCJVw
WMXe2OEPOoUpbcElzSMKtrJnNUXw3+QEnvtPUCUHD0/hwwXbclVfzY9MMmIp9zvCKQi/QfZsWzA2
qbQlPdfnYOAEMRjvfkjbuK/8JW6SE0RomirUfEyTl+i5xIVjWLWRDpcg5QOTjXxrKbNMfgOGPhIZ
rW6/624LTVDl7GpH/N2RveI0N2r1j8c3CEcy7RvykuSPsVqOk7YHQv+iUfmhMsLjjynpTruBDVMh
XAEiE7kOhJFeYKzbLflemCPbAionrTt4l/mFx/GmA11oSOn/UzJD2jvCwNOilgGeBR6YrQUdYQyq
xkqXaMYmh5hACKtKckmXre06v+cmeIi8WJP+Zy8KClh0gfknLG3A6CVmdSR6vkBdNxkdOVZaVG/p
7h8D5gROtvBjhPIIWDpMlgxwBFor9z0vAt2Ki6ugWv4RWayrd4lzvziX2eROt26MK2QefbOF59JH
3JvB+21di0H5rLogInGGzGAmvXwBKv9QKQssvCx2VcmIuOTFdkuqSTq0czX3TOsq5GQQD4t/XrSU
ZLYUjNdmHwWZzHfgCl5xcFM+osTZhB6JNLVqYClvf7E2rPM3CZ70QH4huE8DWFjGYGdre+fMCy6y
8y0FSXrKBK4Vsp6zA9qIl0GuFe5FIxgT7+KOeZG2d4OWT1xGaZR0/nDX/khY64z21QYO1xiiDINV
Gw7th0VRJ3f4K2Q5RmrO13GMRllPcUHfzox6tlPWFWWQ+g5zwJVjDzX6Jg2ffDvI4OMZg+R9LoDL
64a1hdU5dNG3Jm96jY9nJOOnZgNJyYRq9rpZZeZJenbMKYT6iwuQa9nrZlLPyo6AhxPDXJf/SF6Z
syscNRM/H5MqLFJJ7daCBbz050da3fEUnwW5TeOz77ynQVbLvKJOJY4y9G2L5tSgoYDrLp3W5LU1
C2KiSaSTSQzV5SXMQvlfGLlVyhBhzAYDSVcLvHFixLCiE2ImVwmKWqvASnzuEs9wKwAWigQWwRzO
06yLBqLsLF4L+FzNxNEpnKqpXV0LXYn9KWIO/EY5WSNSqOHLcAyJKfwqfWE3Tp50znahhIwch1+E
isS45DwSyoInY1RrAGRNs5o24Px+9giXesas45m5ockKVRQaYuxvqBkuwwPxkVVYws0Icq5NDQWr
RIAMKsXu4I0S/O7hzGbQKaERCBnD87rLCu3UtXcwNyJRsR00hDFEwu5kGKh3KN0DxnJyw7moRyA0
LHOv2gqg2r+xu5RRu2SYuiEcu4AOAHPotae0mOVVEMSGhLJFm69FWqdDUAPyGEWH+xt7NR7X5fw+
rZMr6nO4Gj0ZoICv/jfTh5ZszAR/+GLUAOT1F368qr4N3f9Rl2ExpTuWWmgAQxs1FQko5Hajz0qX
CiB6fI4lGesrRRytPeNAEc1T+TxP8M4kLTxtEKWbpsoc0mnF4cuQU8zOagGGAi55bVqz21prx6//
6gTn1KFE1NmIy+XlmTO8e0d+nthIh1QSnU/nTYYcTvyFCgT8fqBzoB7jwcAuQReSA/Jmw530fRem
LsGslQ6oocLd8l56k8EgBc8B+bb3y9ePmmVbCQz+4MvLifOFj4GgXjSKeJFFDwgUNckWuK79B00E
6Qr0/TwtRfFc2Jtg/h10mCHUK82YhdxxvKtmLEYpjkSHhhRX0JXY9yWaqXKjkIf/2HXSuQ+vbVta
rDa8u3cv+53Cf4OEdO7vsDKHEMaM+EmDt/fYTsYqSPB0NUxrE+jogqT0yakgguM4qVsdZvwX8i+o
TPNrrJJsw/fvOPnhJLx4ZRvfAR+bPEsE72jV/LEKcUQNv6y6R6PFfwPBRfaLHXbI6WloKy1wOuhk
yz+OG+xOk3m1+C7V6udIg5MYN7uMJgRHsEnP9l5Ei3iSBn0uZIvBFH577PWmdgoFGdfPgw1HgSyE
1P3ToQt0jZ2CEmgEBL9hyN2hTPX376s/7jCChBgL9H7SikaIxGVyKnr6KivAi+9asulCypx19dJE
J2ODtPQDVa+0Zt8Ggy2dgexskUtkpGHwxB351OFyfI9xpJJQNl2tNB5L+1eIMDpklyAstMAkGQSb
mBNTFI2UrCVxCcBD6W53dmFeNiO4PLnGiQuPQgo5UwfuHp2lX1N6hYKn8a/yeqMF3fcZwhNgm4zg
3kMkCUxhgTqkbPJozjrn3ikUrp3CACoAbv0X2gXHqGcMlisaBQTvhS7JcokOgk2eXNoi6oa7G02X
cgSks2JGC/F6qLwAWkMA8kZptd1juA9DYXniz+j1eN815jHMDHWefAezgPPMrMr4uB5Q0oTwJ2+N
LMrbpBsg4bxSTSuAquWrk2YBcq4vd6nJZ6ZoFIsIIPgG0x8Om9Ls+tHkZqPJdCrS+II6Dv2ABmBF
AKio63Ie7gTPgW8Tvmw/ZByK1/4ecZ8opwjdhC0GuPU+59MpA3pPRvWEZudpBG2C5bzb037KnZQO
Dsc9jNANIVKK1w2fJSmSZr8oKTJpcHVmquPPR6OBtP2kZ37jFm+hwD+55u9tm7px/sv5FuKfZOJ4
MZZ4oRB+vcP3xwRtzW1L6TPv2ljAT0KXLYwvJWduNM5Ew9E9YKK0HPRdmcLeEgvb6k+OVxms2TYp
UQ6zdntov7HZ68u8hM8UBLDGI7NQzKfqYCFAweDVMJwGcK1ecoMTz2quucTALUIv1z8nHyZ3BESw
JmuQXMq7vgljhqT5eqfx421peEt/VHz68h82N4F4aJUXXkVqLGG8HuP9R+nyBkbZInqpg/oxu1d0
giuQOy0ZOkkMtrPmxHgHHf9gdtvDtb2wQHX4mai1ONplHRPN1iO+w8xvJXITA14ovFS4OLLEyYZC
EbsBWeeNlBEb95QXXD5txc84XFo1H1+ND70vfnczd3FFBg+OKMvWX86gDCNiXQ5Xq2aoDhe0p4fU
7f/xshtQZFeVBbxEY3nonRBy1B3azrgad1z1uPUoNM2dUgg8xx3qdCWxbjgzPSOnIfUupM6SYcLv
t9+1UgEBhI5Fwt0hDB1sGhmK+i+7Qg1dApiADYWe2b9c9GxVnzjvKnyJR8PiuPxzMld54XGo3kFP
XtkQBo5RPK2PmoqRVqp/JZilxawaXrZDqMFNZ3y/8NhRwW984LOIsa/o92Uw5V0I6FZHhZb68rb0
kJ9wpnvLkK0A1BfgCvJiOwrka9AhmPsKW1PYSZKJgYoElbGvOkG/Qi9lOB8wTpkGSOtcVpGCsAvn
bEmhI27DtX4PTJ7NWKxJYgBKllj7w01tMZK2DH9LVzzW0ZYHtFanOWCxLDGHPQ+h2mwGMYFaaPGg
iSv9GbHxVyCpLjaXc5+gXwOPJYMRCn4oc22CBJpwy/G0zN1J329OP3zlYDjLjqp2oN8N0EQNA5DO
1VU4CAwz8k1c9By0jLJrd7JMgeukoXX6crbONnRBrUsQtunP9jKtTqwW/lKCj0dw/J7kf3QUgtdI
T4mX9xTVlQoyoeU1MAXGiepxGQVjtwQeU7Rp/jjTiNtu760aCtqH1+QyiHizTQ0sUj2bWXR0T9C9
1ARV1J7+rsEka1CoowfT/zAqwzXi8zYKcFZbEuNBP83N5pEoEetx0cax6a4Ws+AuSZ4kH+vXOpV5
qwg5tcWHLAAyxP6UcwT4y51tp4DdhYdliiY4BMNXQAFqRtVYLufpT5HsXif5ZE1i+EFEqu3k/TcW
tDj6lRYsyBqvz8frKr2udx5fyTSLHMmTTw8gXSc8kcE0FMJNgSDLwM2NRS6/yg6vm2OHI3lkfKT/
jwovm4abD94xoMBmhsL8Nz926/KndsyrLvCqfLLimo7s0rRAwf01Cg4YQJHwPQVf9wRP53CLRJCy
kS0nuXzTanAx5rIhIcyoZ7m7EV7ixgJSCwO1M6XXfbkAp3xqyTGqn94TVn7k8o2PQpWuKuJ+XbGx
zbpH3r/slhA8YhOiLb7dTDSzI/AcuvHG7fnqiK+lrGj/wfdc3wTzNoEMNo2tExbq9pxGh92y25Tf
dPCCuI3pQFDKlzv5fGZA738kz3d2iNYz1pj5F5rQRjBKHOV2ELOf8i6tj7+vc8LScFakW/6SC8UL
w8plSaXofzyCAXNjXzCrCVlgcl8ynqNu14DZVyHk/OcgBVvkKtSsd0QpnmQnLKbwwtHMYvdRifhn
Md3FY4hpdEYhxZxGvKCscqqb5QqFdSOZ+TYQfuP/J2oqaXHYxqFN1dRrIBLZ6odVSFwkea5/aYvH
LiLNyma+Uxsp0BFjcZjtXT7ixpKMfWOUE+0DOz6aFqBDUgoGgTe1m3BXwVkTmHPxiFzP6W5clRY5
38CoU+FKsUNGaZ4XisP5pybyC4snUDj2NfD9hZCaDbbGxTRBZVx3PEg58TFefeje0ZrMYRa4XzSS
Bh7N+g47C6MvEXqVNZokVosLJYpYHMtpVGlrMaUbvZZK0H4nrX2gdTEZp1ftK8oZk/cW6j0KHIq2
sdP9m1hrbc/6Cf+3+Jixw1Y6olHsSX7WR9Nf+M0Zjkn3OvZmETAzl+T5HxKpMzEClCMsb9v3Pmmz
7ATGtnkV+smRijEf7HvD7vIgTCoAXTO4YhQNkJC2ZBOSepds2VmECZcFtXpLQ6PGLnpaJRXGBRBF
MihLTTFTMgRUccKhi6SOq4tEomO9t8UcKdv2s97C2tR+vccuMAjohc+o/EQtzE2FlFAtQceZXiDQ
SzG91H9JE/w3QPK8mAn/khORRUJHKONJEeTuo3Vy2IsiW0Lij3bKcyR/ENC49yZq8vHHgOPzfqnJ
C73KCTXs5lU9rQtlnINSPNjFYyBlj0qbMB0DAE/LVyZdMoJ2EkBLFhpYekBVo6Xgs+aA8pWLry8J
0VQ8j2Ia0JnokCFQq2n5AAYaKs6NTAAd8RXRkAXclRwnGaBSfZRDp5yiKnUPlHRDBCCL7/T83uA5
h85lanomB6+gXdLmWDv2D4o4AO59J4SJMRWmDrKRvnlZOe9FGDwdDU5IMNyYYVKonQbiiMrqfvNw
4CNA1gqIhf24LWQtQulOjEVi46W3B5gStWIK0rmkKOjqWRHGs03P1NibCGXvod1BG9MaAWLgeW+c
hZjznCiUh/ee1c/H29K9bB/8s1rFr4IEM9As4fbFlevPCoWsq4zGNZbNAjAgr6dZXDGEnrzSvdvV
0IyE5eI/PIJ7AOeEBMjVRIvoyAjRdbMWki8FLxTULRa/0PKzx+eMJsKvz/pjxOSo5Vel8i6hYsIY
S+8F9QgswERr6DrV2CguXTiwGmJVVLLdkZNFVTM4oOkXMpuUxvyCP/A6kn9pZKfTDbv4nGcAKBjv
oTUqyUxw4Mu6uS57Ay32NgzYKBPQMZecdkFEsfNPFMGFma2od7Lwd9KDxmvJ2gh8iRFiQpKtHoIj
oFiFFL01s3vq9eO/fLaKZB7UzobD6+0daNKz6580rzezUhQWeY/BttmiRNi0sWiWbHojKKrFziL2
YKOsurMkdDTv2Bu2nDFosdUUMjIEMhL0X8KpdL8h/IVlFlyQnbnUjnCfUrewj8ESnPacYgZ9/UPo
ayy0EfNM3Y4DV8cKITIMO6vAeujSCv67UR6yydCUg24JlFzuQo3unDMIIBS4bCbRjj0APGA8C3MW
ltaLPXpqUIod4kuHMxy6Dpxo83FVMg1ITgNpRdDkRXriYJnS3F8DO9uQINczmTmcTPlCi8q2VyIG
T8TG80zbzvuJT45X4BXdTiuB2ZNYSY/0RGgpHtsMtdgGX2d/Xc8b8ggSkrtorPj4sSAW51/7tStv
YFg/MmSc4pVA5dnYVBD34kVCE4kSqiCKSoRh85yKr80k9BpEtrmNd04Mm+3W2Tq79zK1NZzgoXt/
LH7YPuYnyl+TWXIH8B1wQa/W849Nfog/kSIQzgBQUC27LXsM8zW64NPEZHQDiPjDLnHAnwp9ecGB
g6cDCutK+7mqpDxNmFkAH7h19TqiAk2B80kheOgiFAskBsu2HG21f1Q+/+AOMcSxNE8RjdNPC5ds
OA3FG+HC917Msp/wsEEFSwHJARfXLfpKau2GU+n3+JebNWK+wpZcAP1xAbf/5azbvpRd55eX+CEo
mSxWhOM9wmaKSze3SacDtqzTY1Vutkb1zrHgcitY0YfeFd+MZOO0b1cQxR/pzI5kqWNsHSo1YTX9
DJarz449gWICEsKNiTkKBwwqNw26sjCSrmxnOP+22OXen09OiHwPXagq/aKV+jPs7DqF8KBzRtwb
JN3qRWMFvS56mZrauqbOq8qxZuVHAr+0L25ReYE+zN7iGTXQnH3nuaL3bvuHQA/mvsAsffaHR5HR
80DNmXXGLAKfk76sHNhofWqnesLMC2YorKyGhaFPe3l0WNzMa2HZbIKKK85Av+8juwlAnZJb/nNj
g/xJVbLM9uUB3ILw8yoy/cX36dXxrvpymMyBnvvQTGV154nE3iAJvKr8ho7/y4lxSHak95KEJmWX
m33no1zjHmmIEPHCaSGJq7FsWSeetK8ZEQ/ERV2oaprRQDgR9Pe/LK/ja+iq4PFLHUyTp0mHAT90
gCuXi6kLJnD62JPJW5Xhx8m2oMiSQsG0V+zKSl1IBxin7nK673NH0BHF0RCqycH/ENhVScjdopxE
j0uvcAVK4WP6z8yXebiOgfhKsrtlBJcMia8dVo6yNx7gSXDMz7jByXvV0REOBTBxXfW2WCTF2c0V
Xe0JwfriKCuzjxKXHLTa7WXq75LddoasckBwu2HvDDbbyUC8eSlsynnw5pF5j/GLub8HdP9F1OnM
BRckH7zwnfPrpvZHI0iKDgu5oweO/c2o1p6Gg4IIGv+AKbVB4oSwLH3n8Ceedok9QxQME6FRHwvx
nofj0PqrfC8v3RttaTXbuIKGMtHw0/jDjqfmgyckyqWABnCvqsaIOrHtSDPmW4lKIPqQOBViLFeM
ztfYcONeMD+A2cfL2O4xCxV3wWsGc18gUKtqm85l6BhAwlcD1qhKHR35bVEBRvFIDfg5B/Ql4HVb
GryN5T6TTVQSBmQRG5I+rbK4qGZTvTSb3SasRJ2D7fAgmdyVM/ohJhRyEpJ4DiFgdp5O5tR++ETo
7eTFqw1VyNTrn6jD491sLj2XBbNWpfvsDzIRR4vqHWC2PWFTykfhm7o/gvNbazATZQpMpnTNU1t1
XtIDLFCWhtGvNLC/Z0ltdPFFcr78R2d0LvjzSBjwuRiJFnPiFBghsHEhGXgvw22V4/flSiXUZZpL
6sslVdNGFE0Qrg61L2hkLDrWBwG3YFMe1i1KjuRnKjwRglwb6XVyem4x8XWYryADTvXPRyuY16Re
e2fePXby+WUR3c2D64VO4PbxXgJTsdNvYGznXT7j5GdBfk/fxsT+E09UQske5cWGRSe6/M1rByMW
I7cZgrCPh05OUSnMj6xgDcqSpHHR/cJb928DQTTtzjRUJyNWywk0NObTgOvLmZx/D4CRD/0OE8Ux
ADj3obioff7HpisfFArAflc202QUUTgBATRp7YMmWIz9/0AuBDdbejdhxpo9bb8UISv9Y9BnMIkL
dC3zUJiDpJKR9Lk/tdQ2VFnc24lKigtBFHsYKeJasU28F3KxBNpZMQVUrfVFjZyxaYEMtvAmmdO0
GnTmbzxRRSntyD12Fd5w6Q+OZ2oXitzaq/cu8ctFfI4dfL4kBdCw5dOfku6rW/h86Tl7wNsNIrW3
Fh1iJ2r6WvXcVTsGTp7T92wOWXZQYUWNDOjTTJGkN7TMCq5gQ/ET9T5ZQGgao5zfw3XOHDG8pl8+
bMxC/Vgrqy8yZKTDNbN8vmJYTxZS9254tisWoZP1WeOjrN+FmdSBH7APdX1DafwZT271+EoBzXg8
ae5S7N28eNM0T4y+V5UK46nFyIQqDtWT7kE/Zf9+v/I3bT72GwgPmp1/OfKs7KP2v3xgfXIYvYtz
3DnHWf945KMsnOKyK/D1VhYyklI4jaT/ZhQtVRtPES3bdCLhOWv9lE9psaYuDg/xESkg2hvHRKl2
M2lJCyumtR02SInQ7hv6xF7RCVdjUShdEyq77dyBAUwiJIbQ2o2ajAtvr7YBOBCwY292NTPVvAtj
62ME83oduxEqWV2fozcvWYiKNFqcY+Ssiw+QhCDnkBLtyGaW22lGHe8x7Z28fvqdxuxiS7SxYLLR
mwFjguU/DdojcN2mbjDLtw7B+EygDKIMnlDVSKwRHDL4JSgdduvtaySj0Xz309X9C19jA5SB8+Oa
SDuFE1TZDnPDW+tJkJn7IprYYkXvZrkGmkPeXH/7zo0lBox5fTwqc7PnFebdf3IJSkhRPr6ql6Vf
I1+StO4EzQvCJyj8VKys/xe3F3MQ9PfIKxYm/g9Om2YZCJ/pSHmkhp4eWmow/WX9Yy8jhoNSHPAO
pJxPB8bk439Bek3GpfVTtzLGPU8k2MkfbPTvYu7Wak/9p987axc70T9HNac1t+TDWTQReJbd7zbg
w8F3lFFsU80HvvtLSBpObI+XD1p37VDLI2g2bfsRhyHB8tvlti9hN/QPOhRDI8HoaBWy7CHnV+Ub
x0rJaPRz4WsVGzppikg7RljUh4+qy2Ir0TiaCCM/JT2W9BGeWkiUcw2/mIqaBpaHhU176W1IHKVN
QpJHXWgoexpqwJ7hSqrMWm1/T9UwU5/2TJZQGdfk6SxRcFpt4mCusKg7zLpMp156NLF3sYJ3x9je
tYo1P6YCKR8N4yQEmn+2yKm8ILAkNCd6skHThqWIw36ppesA+LSygMsmrfqy9+YcfixcGT+1E1jx
DUD7ctBx7W3BOGv3U2O0WfnJHl0vRv9eveUAkrLYX4zg6sAJTXrVPntgKZpmV+s1S/lBeOJWVk9c
VugCnkQb4A/C9zk7Sc7KZ1JFq+DTc+HFrUtCyTXTUIIsSCOoaMfg4WmTJo5wtztsV+xj49nimRaJ
eqGTquuQ+CI+H0672NyfmtfUk3kulWIWwL+vJtbJnQo/I2nJsBvLgDUqNdFuE2Dsq2Mu44GTTqsB
OkeSV+DKwRyZFzp5UIGv8Kl7YfYo7adRIRcXx1bxFx+y9XRfn+8NbJZkHWafZOXON7J7To9gfQk9
xg27ZRhHxp7jWRzIytzSSKJ2mWPdHcq8Y2edFOPRT4crSrvQU3us/0pudh3iZ2VGtUtquViu/nwB
JD2yKZuDobMAaDoaiINYum5x9oe4TGnOcOFlbDEhh74WPBv2Plh8tvi+VXmfswgYUHDLqdpINASy
ftI/2V8CzKerRtkzpPdf9WpPnUeyKyfcT8aBnSgzCEmB6iQa9mN2/aTtnfk1ptQcFukamkIsAFgp
YHcPL6pPhdZl4IYnq+3rqNwnInmJhl2821kIZhx4c3ReXFq3RDeLoXHdTcvPumRuuKJ+CUMM+JoG
uZdEDAxMS6rUHOl5wPuI367EBswjEvSKcmO4muUegEZM1Pv07SXjnRDKMCk3OAkS0YEIU1n3leLH
we8zw3Dzf7t/t5ubxcBHcpw//hkmQyYggkeBioN5S794SZbbsiA1WxGnZoMR0Y3xHbhQuaaKxuoh
E1kn2tl66NHCvpCRFoAENIER4KOseGaJHhrvRnzCEkSY4IXVfIOQ5m+KH5P89AuR/AFR2YocxiF5
FIVupxRke/V56x7GQ6v7em5t3AFCvlZMfG6emaHOB39bLYjI3AwyWVJ+rOIG7NESMen1uNmjuz7O
WM5Mc9S8PX8EpBoIQQkeOvf6S+Bp+ClrNBbNVZIRjaMqJjUpk1MMb/ECJF/i6Uy4uGS79dTm2zjy
sS+3EFFhnDlsXeDPmGBPWdl40JKW4/5dTCKPND/vYTTE7+hLOMDQ8MfvdKLyv3bzdLGCb2NDe62y
BP4hdaDBj6z1nELYGfoKiyognJDoBhPwv9rgbmwtqgnzlnC4/0DQ5keu7VR06kJFDckZ/79xBZV6
QUCgAqm5jufNhgK3g9P4+B6w2Pt5nrXNbEyAfCeJaewv7K+tUwCu/zSy62LqBb9vqCWR8cXK6H+N
hm+GsdLy5Ns7gDg994OAvgfKGQqB5aXcbkRUVQCbWi57XnJKYQtvVGHdiTfi0mkWYZKcyiuqnWL7
fW8mL8B8HLI2Q+XQcJU2UJdef5teIOf2J79Rfd3r4IHYLoxpA0gDp5AJbdE+VW0MVmuHzmETl1BP
XaztGMIsXrNUDZvDqfrCT+rq6zxRXVVRLPIEYRxxhyG53/+fmtZsJHOvh2OgwhGRocJv+T69rYfw
ORty6XDq/DTjvFKvq4t5mKX7VOPDyRECjm2bhR2z8YlroHluYNNxqthUuW7w1eSN6CUZm6WH5zam
lpcqcmYf56NZ+8UT9V20ylsO6i3JusmCBTir7EWY0nZ0u2jSrihB+3oBSPtcxqVbRBUMzMwTvhdY
dsqIfjqK4Hf/S+U9AlhxrEhTe7epJ9s204aajvBT/ujmy6zdR5lCh47hkj7S47U87F1jG1nb4ixI
wvmYCVfdgYWcffjB9/3DfXJFwezL1rbzIDj8S4aA6J1XwipqiGb+ECxPp+XrYn73LeyfME2zB6tv
a4J36ViiVTJweEhasolzilAUB+1Vn47wgkFeN+4+FHBxygMDrKbofdG28k86K7wlu50d0zHqnICS
7ZDxMK2YAR4DMkNvTW8Tpag0/Rp+AMhnGw4n5ZRKIAQIuvf+NLQ0HalkbVKMZnDJajbWEg3+Ay0X
yG8TRI5V++Vx61y1CrRcHfd9RcDMA6NyKV1LA5awpIshgP+v7w6ju3ACdAHEVOFElZcG2DRsOkJG
s7jt4Gu5WWb+r88zhZJjU+EVe1vOINexnHsval2A0GCR57bRo1mr1+Y+a1rkTjX6uJF96UiFOfPh
hucwZrKmlCgPfzcsWr3/yAibOjP8XnyLIH8wtQGVKZb8QjUQZs3O/nj5+uN+CKzTduqdAgtXG6AD
MDdwDdsE0W0FLkE5ldQOZaoDl8VvUtJUnnBea0Bw+qG+KGmHVVZblnvAQLIXYakUpZmQiEiv3jjt
grX6jKmbGY5DVU0GMhdzOj6+F6I3VYq2rwbIxxC75a0v/ZMCQUNBZ2qKcF28d/smhBs9bGNr0Vne
jHzvV7R6OWZvm4Qi4LPL/nVKMAIj6oh9t4GzKSiWcTPBH4whoqrZdKfJUJD4lQNY1Giq2GE7uP6h
+btsFjdpDMj6RgELMkLqop63cdbAmxeGUrYEMkuIIDs762bv7IoWdB5iEWFrDAK9zvNjAplP6Z5Z
gvLlzRTUrfMhuj5lmNF5BtZJXLJoIFx0+TFHZ7JLkaFem3FRGoHZK5NDyLzE293l4UYUGiLs40DY
ZVqwsSw2lhuZnUYrrblcgS8Jrtd0utG1E6Vrfji4bM5aR+mzfhUz14bAqHJJXlECOPaAqUmebkhW
tAnLvWsk020j13JbhhgnVmCBgWsGYzOTeCqR49Z85WWROk/6G1PYI/+bIXksE/g5DIcExpCnEhPU
5RdRZaH5bbHDMneEuSWf7OUWfi+y1RmRluX7X9FJr+nVCBoZooaIxl0mnvpO8H6ejcLbb4C4CU0B
fiz3c41RCY2Ckl4adW2t02O35yuDpixJGq3JVmTTo2w+ITIbxA0fyt9co3kc1gipBwofWhrQ4Yiw
P5DWTmSlTBJTaa8Gh4N9x48B9zolvhJkYzHep0av1hiZFw3r3SrD31CHOKg9E5n6XxkGpa5TJcil
15vGYRJUl8XK4da8RTgjxYc5MrDRGGoHLI6kVQZoL8GdAVngjHbrUHhqnjzl3Xw4G5SYDtAEg4XU
zoM764J2rYdkZuSsA5NP01AgqlQnKtFF3YhMcGbeEC0biIJzoc5GAB+IrSw6MaX2aDn7rp97a5SW
JQy9i2w0hPSUmSCu60cwGliNe8kK2J8BQePQBzcK5wVi7+f+CJ8CC3Vx+BEH4ZInsEoQRUMsRWa1
PJumx8MfkOCO5ONM9dazMIA47SlBshxHGTPBDHgNqKnRp+DsUQIksyCRcpiinEtaFDchZrUokxxJ
ZEZq5R7yOLC7xDHtY3ZAPxVN9bJcJCShgAGWVRkhoTnLrBg9eZFWB7O6UbA5jEk41Jv+QgWyc6mj
DvbkUHqPTITKT/xNEVqyW1NjkfQ9R1gH7cwc8PD+RSYnCg8eLu0Z8hp5Jv2HTzUEImbaoleaN5ho
MSCQxrT+p073o3DLTQz8NqpSkw2oOKMW9ARC9XLpWAk7/UInfEulnIUrZcvRt7w24kKAL2HKC8hT
uRASBxgGTQ0Ey460TUsG7eO4xV/PQucBvtp2UGsxcmGd9thIWFYOir3bX4mSVW0tq/wfbk1l/YuS
I6nAR3sTP7a3S9hVjGrGA7Y5KXw8eT3Oy+7ezYLI7DUUmMSq0jD/J8GcuIK/6wI1ULL6vejdJ5am
xUY1/ToyXk1GGTi6xjkR0MbxPCyYLrza3CBuMx0rgLaIaST86NsTQgFYrp9noIK8MxF+DGio1Vla
Qym4E/Cv2Rp4rjES6GrNsQ3bCXgilK76Dnf1zyTrkErDmlksT80uddtQU5kHltE/Zaa2Gm2X7tXI
USVDxW3FLnBT1/EEUsJ0VHOyqdUYbhBrWfNw46wqgxdzPePCw6s2uHECXD3teg53DfZ+IOkrcOKy
czgkc+p2HdIMN9QkfuWDJBsP4law4ZEjdKjTpom0w+SxqAj9SU64BkRwGII7jykt9J9tTIawlkMv
u3JiXYmQFmLAd+wtOtzMkIqVN691qi4zkHO31iZOlv1uCmjoSu1BTBaFuZGGMWcUm9WOtpQeH/da
uHJdlJdaaD/L+6AP8f/5mUL0rOTdvBPSuWp2s8Is6RzyVRYplX6T7/7amo9jUwXM5p/gVV+2wBsf
J1k38cYZYKFyj6Rzow+MZvDWX/8qzwkXgBkkzCymQr0hkZ7yWy2Mcy62fJDLbX7ygpNUl+S1X8D5
0qZLwzF5CHJXxErSfeTdXHFkk06dYRBttbzciAzK9PgLvTKFrM0Tl8KZUSij9XdugPx35msbRorn
XuEJvTToB5bjb/Icpo/P2/0gwp7Uu6ZUOe9KpqrbrC8RErYNInvcXhaX2abaPV3UJ6BYDkaFqcMh
3hqnB9jc8ig9C87esIlhRzMEitajzm+xOOwFIIcv01xVtCK0f9WJQMYMnR1+xBgMnmv0jyg5gtCb
5JdPenG/cjlR3W2sibO1H3VpCbWamO7JsFIMDLS7SYTXOBwt5/3csdGDj/r2Rpyj532nuos/NSKx
oBzZ1ybEoE6PXgX9XZ2PJep6fSh22k4/wVm06MA8+QeXzGmUicUP4BLZ9qfbpzC1tExPG5uulRDQ
5LALWDu0Jz9O9+mvwcXrObNmreJ1z0kPkm317+OvOeV+dZy10+RRhOprCfEgIEsMTJE8DWbhSHF0
8nD7grX8+3LVoNY1KKZbosUBUTmPOrsMe+GZTyOuR9D2ubG8Kkh+84Kqr0SD8W2nMKixfQuG9oaH
uvIDaycYAxo8ldCOtFUAgYBlFrWxDDbarnk7XSvoR/8nrFBVQ0rS4R5j/7g1sEUJOvN2uoN0bwZV
ygaueWSEQ+d5S+w/H0Eyj5o4JwtP37GtluHu5uG72vImpNok2hIL4EGF70uI21HC9eM6Avlx0gI6
L63wEfzZPBGxFCpYNtMkcXgSy6HETfdFcanYl2cVtq9ZK0YznzsionLvPZiVs7DHoDCsKpTE1+Cr
UYfcL//+8AdMIBgN42K85WPiUDZdz9r/Eezqlt+TCuD8UOlTIgk5xHZxRCYm/WZNsQ4V77IidG6t
P6DmRfPDj3tPeekc25NMF6/GK91uvlH/cM2Z+5cs3dC6f9hV2VSa0eq1pimjUUnoPY52JqD2bJme
q5Ff3oXsSiVi+Zpnn3ytRyX8T+0ZjeoUrTDnrJ1KTvrNuqsBemhnOhCAJG+Cd197C4k5JTLeHbWl
5kLX/IiHVMGEYYHrzVl4IMeVxOZYHAQu7GsobjldboNBQzrzSYAguEcMUZHt8owa9Gmxe/ttIk95
9gmZJKl/dfMEDJQgbHMFteNVwRu1gU22BFoKsEq9FXdhmgfJpl/FMQjUyMLaY+E4JiLAIhHVamdu
wbYakULVByGQtHw1Xp//vph1SiUfSJGQrmBRa8deM/Frddo4qG2cC1bc5/LxuW1PUSDPAgrV5128
48e29lMdEQ8CC5Lgxbb/pmxPsM5pvZUxCixtb219L7SsCu74bCSdCr7FOF2c2wZU9SVN6d2up8RN
P8dfxRVqkmL57BylTQxBEBrkIY4/1RxIMX0cmKKc3rSouCg1kMLv5lyvd07sIX0aw8LILvYf0oCa
Iyv79xM/q1qW2KpozgAcc/L7XdabkWLN5R2dqC6sLyrKBtPKlD11JgXhA4xpcFO5aHi9yJEa6/j1
txCcNq+OuaQPfucclaQuNwPlJnji4N+efdAeIbM/eE8QyH+6IvWRwhssTf3ql4PLd2hfxsT3FAo3
wWl7b3XD5nVtDZ8vog7Gc7cBZANKQOVpksaVegkmyPMQSmjfQrcXOYKQ6MJHvh/S1M7hjkyS2IlG
378dx3KWB/6J5osiStjscuVd8/5XmX2Y4utxx0BTo5QaS1fmXs2ve/+Ufa9BaGjACvrdGhuVdvrd
DHCbgWXInnKYro7RIyycOkO6KR1phW69oM+27xo6zqHxt53wA2PJK0wOwiubbqxzl08irUDEAL9z
4PXkrnW+ZgxhRMpwPn59fxmn5UZ+0RbMoFs9t09uK4zY1MpI9E1y9zl0psYXyaVLzbmq1SWlDHfZ
H0e/zlQKI3plMUAIUIBThrSrmAjwnpjYd0Gjzoz9nl58wbDX4Ynd6/cJjjpfrIfeAsGpy5zCUpVF
fp8ND0rYAttUSkHs5Lt9CaW5tvc+AIubsQO500N84n+4cUzXeZeWUW+yDd8TQKJ8Nm9Zbf0D9hoQ
7Tfe4nVycNwF+eaZUPiijEI758qMuw/WyGZUxRP4sWivQoHBsQzlSkjShxV9wJ7Jlsek2yaacNm5
4ctHRdRv1A17es18LiDKzzhHd5Pmolg2qIT/GFHrrPRjLDSdnfwgddWjxAaqcr+jJ7oANSVhECjQ
qSeP152nDsnmwEiY1z1f1JvKB1UyMqLcSiK6dVqHK5m8/Wy9jM2/0k0Naa4VGxNySrRdHA53q+Ma
P21g7IXRNl9yF3PiZRyumFwyUEFyn3qZPBVH7prSFdQ4R0VLKgcde/STyx5g3Ppy6g+ZeJZjD+DV
VcHycRtCzbLo7kLcq7UTxSk/EKmz/kDMtyQAbGZED24PIOSAj73ZAjTEYTD5/NpVn/fSyP7e8AdI
omAR6MLj2omVRe0j/Vkg6SKXLp1w8q0bMaYTHFQJMSLRef1lRkP/odkjQFHDd2z8SyJAZaHTOmMI
gV7u8x5XF5GCd26gHcXukZH8XFLLlpRGlxnxAYk85CMEJyLAyigmuOCsXqGO0i2h0LaWM7vB4vbl
t83fkKw8UJojoJbsHwnJ7uxoTdF6Ncw02bUphgLJZCfHCG83SlLpq/SjretTWlamdpDg2PchchFB
gis7uWx9O9guIu1jtb8gHw/FEBUq1+jw0qL+RI9QzNcMFVprFxF7aulMp5tWqO0U/hW7xcJzv4P3
b2yVmlcZQ0SXEbgr/+jGgs7gju4F3UR/nCr9jx8dwWcKnO3zb2k1nKtf0ZSIpHFd/nfPg27Djgn3
6GgIRlJGvwYYnhDZOvldvpONHykNOBPBW+cNonSCmZ5XRs4M4bl+BxPgU99bLUaWO0cSMVi7OmHk
T4oY6eRsGIwXHZZSIh+M0Pd0+V43ZJfFS7XjDrETKjDuczNrV9rw9oLZKqMEsno4aQfOgjPLjyBV
H1N/yT2Wy9Nantr/ZCXx3w9C6YXw9JNo+M7XMUnZHSFNDCN9QGbh684IKtd+cssaH4MU025fET0V
5mFtCfTfYLK8UV60heGTfgibARfEiVwV9Wfi7w4W0R6NYfHDnU1x3+Tscl9/5UTFV2bcXa+nIvbM
L7rGCbiMxtjFX/OTsuPl361rp7gMjCKaKmLZkRoigQ+PVcMLDgfm/mzTgPX91lNGn/I0E1+zxcY7
avazcfBc1s6SllZXwx6aKSslt1op00Z1nsnYzadt/W05e8iwYXjHf5WZTEx8lhHlhDNV7osvtNQW
HuReShMAfIRKPwRhM/iNAd3+0WgDmUrtGfZ74KPtzif+q3UU61rvDIr/5ZheQtyuFe5mk9NmMy7O
qiFP4jWqaeIYtBl8klhmOneN3zJ2tKHnjBeK6u1UPtZeWZ0s1HJyRrtSuR662MQLrXi4NUJBIhbP
PyS9uP9k64E6gvsZiqRt2F7v/1u+h05nQA0JI6BlcGPw3yWiN76VQOUi6oX6TtooxlKU+CR4SdtV
Z30bEoH7bPmEnLj5BlPtf419FdlGRtXKQxhW/1qkGbUek8yoAeLfDHNcuzoJmQtCRbDnAvKvmhvp
KzWzmO7l6RDwAy+d8BBBwhf4kCmKG3pCSh41WPhLfMgN+pkeGQ7UR8aQb47SuGOzhKR93DoFA5W8
Yinrlcbe7uPwos3/WOJ8003UkN23eyYBdkOskWB+TRocoImH3t3U2aXn6s3Swx/jsV6zjTC/MVHR
xgn2UNOx53sFe12UUysqF++iIUIm/wwOt9iMMeQjOkxafAHIiGSYuFp9AmrIqTYrLX4JCIlU4xu3
sGZQCvw10nmm0G+nSTOg1w2lXZ02AD3OZJFxKV89WOPYsyQrleB76ykGJcnURiJEnNrK36eFlsIn
90wu55HZ8h8QJTAy9dyb59frs+NhqpozOcp/7EZs3ju7YHb5epq1aj+qOG8txl05stncjXIQdqI0
0EJxEVbSCpOl2F3itcBBisB9bp8KqKL+YqO8ApYa0zj6P7+qREpHe+LQQfCuwqJ7/qqbzLMzsJsl
rIJ6y9Nmv4R+bQXBRjds65eyxPyOyc7ihi//f30lGYPr3wbMp+gqahEhFegaKEHq+JVkW9Myfai6
Aep6JQuWGDx+6so+A3HFyW14gaBR7DhV32PcmhnJCDpd3YvWKW34kCZ6RPOTQTPfqWWTt/g/HazA
L2uoRAGdagxkyND/QgH5RLW3Lg72bOinyYhJL8bb0Wj/WjagNGU5w3qCAPy52CzGFFCVMQ/0YPrk
yh/mvXgSoBZZU+wytY5gnm48O/6rWG8Kf5a8hRSuoJ4FRlqOdNvOVOS6nX91LjUdd/Qh6wjRQ/g5
8gNzL2mQY9wtrxc6b84Q6RQwTMXXFJSzrjNbFW3K+fyUzeCayTKqG6P3pxu+Fsi2g72KLiSeNbKE
AwD4yC4kcSRJ5VJ6Oi0KbdqZgR82kbMVQJk2NXo2zk1Y28oSXdl3Sd6zXsGGH1o3w0CxmDm20ROR
P6aJ1bTdWX/OBYLWqOQVlCcs4b1vOjDJycV1jqj7ZYK9lMgYhm2+twgmMf/EN1KYKpT3FRMtvjoX
WhXBz4ky8dNMZCmC5jEWO5P3L6T9vF5Ogogsc3MSvN0vhW3iIS1oXnpFgwKmdVw7UIAvZdr2XE7R
gxMpF+8PJdek0I8VdTk0vBm4AnLxdEd98ZMYywmAvl6gVsGv4rGoXUG68gMzEUcUXvhXGBZZKPRP
1B/e9BX7Yw8EQSY1bWNnK2GvxBncpUnbAdt19DPKGIRYTcXZN0put5P4ObHBBQ0gMbJQ5R9fryK9
yKLhLC0uhK8KxZlL26AQcvtsRZEGVraTBVYYH6ULfcsFpJLHZOci3kOX5IUcZWuqb7USTl6KWmar
h09LDLcLFVmmX+M5lcUItOdXVmClizwm99Nc0Qd4EzHjYOFYcXypfZwY+jzRpf4Svlgb8Su7f5b2
rV9vjAlSH/4OqfescuOnR53IO5WHC/mEVrfTP6ar2KG/eQ7ErRqoPR1OEiJGA7aT6gyioNtZnLSN
7f2QJn9L2Um/lVeUjnJWCsZ3qnGFEQDmd5Gwy957H82AziXtSV0xxlETBoxIFXEVlgYnleN2ORKu
/A1tjKVtcZ837Nkawb2lPlGCmrStVr76gk0BXviI80zgv03tJ1WEazc0cUczVZBG3WBRTe3ohqTt
V9siac5ndXWsQe9tlWHbv/pZGol1OwU4t3Ycsgvs+CWbS3QxyU8BDnvcXZMQNcsakYApaI89eCeg
PUDIVAIyEvLt5vjrd4fl6t5MD2x+l9+l4RJqfi0a2EnlNW55VBFtsqs0L/M0Zw4cv8AVYOOD259k
XfL8wF9itrBRFUJGcTiXRefIFZWNKg1FxmfXLBoPdm1DNjSi4LSYeGrix+YcGq3Jmlo4Zo/qK7AN
nyqnuGSCP8tT17pnHGxbM7oTb3Kg0Sx/4WEDNkg9Ri8cS5+XJ2lBrhM66gFO6cnXrYV5+3+1ps+G
h14eDh1S0sXSQzuHvsd+hM40Q/bwIAvuteCdlRY6iqgOxj0YwYeNmDq1CZNPtApjc66f6tKaU0VA
p6hpO7JINJn8Iy4Qjuv1oSKNv4isY0TUpiaqT7vKfuvjEWqG6Sd1/W8Hyw+RHZb4w3W1V11ifU+e
rQaQ/M20oj2ixASZOM301CSKYbmsLu/T1WDnQRcXeX0EAudjNbMzV+PjbBIclnv4Khrb29OWTreS
E07p1zyNe1EHtBgqIimjJBt6o/lCzk/Jy/ba7dvbElYX1Fe6TSfjBQCBBf++hN2Lf3ErIdPG6ALV
X+7QlCr8OFRk5R+cO7Kbze6d4G1A/gVmJyUn8Zm0S+twn0YgyCxhncVyQ9toV90fBFCCwgwb+DGs
JchnSzPewwvtawCPMPwwLt/IHs/EOKQwhOHCg62KhBLCqpO1IiPModykzxBsdb667sFCkjN30d50
SE/Bm81D3EC380zwxzSttXAYXww+nxai4J9iKhh8kvXNszu6mK8Dl9+Ki6vfcYOH3gsuQOg+8ITc
K3QzJEBvHDYpPvb95QZGGRqU5S9Zu3nk6M0Xe+BTZ/LV28jM08/ORV/MrXtW0RlzxZwFMkfXnNZ8
F1n2mWmXk2WizjtHPz1e8VGXvHEvTKTZq3oQIwNytAUGFn5H2oaPLKbLDCHGTe349Dc2b3cYLeu+
Bey9JvO8Z6XkbsmtZPV6wyrsW1Anv3pFsnxPQ0cWxVE/j6HQ7WIfzx9VWbqidwViPaYyUbmDOJnW
fh11BNmlbMSWg8l5IZtIedukFV36aWwtWGO5FglgCabS/c98vzsTj2WdONlifAfakUj2mZEFWJbZ
VIZ4Eyh4aI2xNPG+HYIY4PDQ4p1V2GaPoYKKiXhIWEzGXw8VD34gHHj2NZ+Zo/nNL0yhoLmLfSkv
CkMTKu7bEetfKUIXce0Y897GfEycvfqYVWsVi5eDwfpR1IgPA+y1umpNyJsewnYBtFrFenKmSlLE
ucGUVtKdjWuFxUkLKSyMKZJo5B6JkYbyaFA3QQNaJ3Rq60GOXqDVGYOayT8BUUYD/T8Kgokr5BWX
ExzJ9H+AHSWDJ7tg09e8RvSCBsErU5/H35ooQ4YW4T1s8tJlDWoB7X/M4sEftWBM1hnfU+8nHGZD
23kMPV4sg6lNQcBehqrcLRUR/tIUAuYg/oCVjORSWDEVJYY9/BKzO78h61uudc67jv6LRgDe+cdN
7aQMzhKyJhkJukzGL3rlYfYEH7TeRcKkjWGziK2DoaGzEpheNNAuAYAyYZjPeuemDz5UCqhqyY7O
H2r9MSdfgoXnQMxOUoo+jz6D0ngXDbM3fg+N3Rgqky5Ro3ZXS9QA95CZIoXIj5v7INba4gSAAg/6
D8UE0BgWZClaDCipFdbCawxOautpVAR7AiSkMVi5hhpDZsAGJj4YIQjyCLlA0TKreQ0VV2BX33sg
YT0YC52dIkA/9uo1d0v8ucAZ/pPxtaTB2WUOJfl0sqXklKlpdM8pW/qLUN7Y3nNGeWL7sA7Gv0Ao
FzgnTOWQZOQV6PulErByIkaAED3ksQKt/WyBLBVsg4o+aANnbImgZllwVtNvs1UB/TCoIjebzogu
upfeX01pNW+nxQPGlvN0saybqOqZhSOungMtXPRqsEy4vs1S54E+mAspjLrEtBPTdZE6DCB2DYF8
OJbwOaoEElO9ixg+fw9r9kBd35eLIOdvSE3086bekGKEUYNz2uuRZcLOdscNtwkrxOx0cjwL3US4
yNE23cqo9GE1EOToqpYWGXT2Xf6SyN59c4oWWvekydJUfu65XkkRrjB0MUzHGvIMrw45Mu+mHAa5
aUDrEJ1rrCdLM9F1IKkYRx9zd5Iii8Zau7L4XbX9Al264NDNpvqrya3s2nJLlVrr6vJ+1rP7aWTX
dt9N3H8eGmW+kfiSWC9O+Bimo5U1S8rcup2EzXYX9vTGoUfytb+xdoEP6KnM0Ii5WKJkQwJVU50a
eaNgnQTKIPS53RTPYOOF01Kyk1zc4VpIRnRUQtaaGYu7I1IgV4MbeFqsOQWdL88gZOJfxctBrqe2
ZZFMJjQ7X2r/OmU5HtFRcLzkEiDgFTGyF8Zav7lTCngkVSEHdYZ0S1C4s7RiZPUrMM+eZJ8p3/Kh
jjXLUF4L07thZGaZav2wtco1G7EkNhbnUKGts/GuaGxkwIZ9eBOfVIFn7USpJIaAxQgD8h5VFBwB
ddUoGCBKqWwSvh+Gww/svhyR0WVVMicA5pRB3xffcgYyl7sXKMpTCh03K9xmldvQVPlTk19SrO8d
b9EHfHt4HRboJH9jBovz37ATHcf3pnKYswQOO97xZ6ZfMuK1+sSy6Y5+Mnkz/hfT+Q4q+1AbbrIU
RU/btJgX46s0ZAzJ71djQzgxTCp1UrdyAb5xJk84WwTAJi1hBBsRz8G9sNkjOKv3dooad69/qma0
Drs4rvUlhyUWHTN3FOD6FCDA7wVMyOsPeaNP5jNgvk0JWZzbhD7QPr3Bw7OzqI36gPG88PiqAKAj
ptU+uJteXRnIIA+yRKGgfbwEdHO/iDWttg2LoLYAjG2x8poaUTOBu2/dxygEUTfUFpUhuOwJ6P0a
HCX9cqXjxxcfcoxbd0p2CFCtZizYNRW/IGjH+8GI8xQsCssotbA1ep4391FDKRsBNMhpVYUuHdr9
rxtucuR6bUoNsyvUbPKj12wGyvasWojnMpl1G4Xz4YU9v33XiWuiwFMSi3Uv0CXxsFBU7NSFSGHK
GJ2UKWj3tRCCzOUQSeijbW3WudzVR1DKPh2acMxyePUFmFst44edzM2ulDKnlPjJvOD/Ai0MIF0o
cohf3x94Rw9U1h6CsP+4qFsjc8PBwv1E+4KTJ/xgDC00C2yUAe8oPZGgPTws/mcpdmfgRK/SstJ6
/QkMWuVnf4FrcZE/BHjxh4lu6t64jKo9LmcBua54Pr6azKcMsDlteI6634YZMrmtth+0IY9hQuc0
FA30DB2C/ABB9lGfkY+YzBhy6l0sI7DJQCrbNUHsUz9O69+ZHOFR65f1P0pyoFn0Rnm34/2mza7V
II79A1Dky3SRX8E8MkSRliImeVHu6PdL+olMLb99G6aJM9RbWb3/LJ68jaSLYRa8xDxzeFeTPbW4
VQrbLceyHf71gV1jt+99Hqn7lV3J7hcYbKdWwypfS2+4euc896aCqFuSi5dAbqSU9HIzuExHvvX5
QzIokZ8pZYMNkxMEbu6CRaSLbNBze2L/e6WrD9IP8kdQ24AVcXXHgjT8h3R3j5o+gB46NFiGev8N
zL6KKvhaHPOlJ2KUkRifLCcve4XvPIIl5Biq1mH7cgktRUE5OFJsGXjzGS5fbZNi+PNczdNEN8yD
rnIY5BbEEpXuZzLHWvgeU77mD0cGZdybaBKR0cu663CMNGdA+nUTj1LokxDMsKBFEYqoYJidQQ+6
OAent3cOr2DSH0y1rNyAVPeNXyjr0CX4R8RXoqHO208e4kB+8vS8pE6B+0C4gAFPwCKmslTL9Dp8
J246xgT+NIZZbkWrS7E3t2eVEeMZVGc2CjE4t7eG64k+msW2RvD1rx7gfy6RsHmClva2ME2YuOC9
l4y2nIdWDqJVJErxymdAJN4nsLSnq8QDY06LFUCv+aLvLYnclImofUDS6PMsc1Ukuc6JUplPdg75
Sz5QFNAxpUmjuk/PiIpPGwrOyRPtNR9jK9f2Ktp4dnvkqR8yls0v2OlRELJr/U1r+hERGV5Xtkuh
RLfQ06FZw8XDswXAzvblUKLH/8QoSiaix0FO63NSafBJn2GDrwyUyp4uySOFqbT8HjlL9mNOi1HT
XYgDrwAT/a2S5Rs6Ws/moBVGj0SrD5B6SGyqdfApGXGkuWVQqEpPbemkLh6bw14EudJThtlzl1EQ
bONIQEZJVvAm2amMETGimA7G3TyyRiLuvqNY7yMJPLoU2syK5NWR6x2awyVZlmnnEUrhodnUDlv3
z9k0JbrWHP/j+6jXoyKM8pR1uGAfQUvTZpYUyMYCnp/Ltu8eyRqYin8JErsKg7vBhShAN44Bp2FW
QI9kYKAkLqm9k3fB5mcrryODTPL6zE9EDF6neC1cTOjCtSpTcQ53eAAoe8fP+OLZXLawqMc6IFWN
Vl8wsmFfzI0qANXWF0EtOynPgxZ/Qc80SWxokZ0hVzW7R7FnLhcIc0QewkK828yXeR+ZIn/N3Y0W
u3HQd8RmnQP+JBz/xRbvRN/io/AeYyKnmHkvtSYzAhv6d9JDxpbQR1txAn22ys/IbfJAq5rbnQhQ
TdSaeeegygknUKGh7fLg5hjwjaIPhqBGzJ4KuL3QJc+cQKYCn6o009I8JF/VhWlmwuPyfopJ1+bt
9rhHLKg9ui5sQQPJRTfE3QsbOVsqnnFvV9eeLhA6G6j/fRrgV8sM5mqwDvngI1f3fRmxG5CZkGdf
okAlehjLJThFpqS9i0uqFVyEYz/ZBnZm7auUm+4Agd4AQ1y61i/tXsFvA/hsJtbxaTGvlahDt9x9
zZ5IZycScsr1AmOQB2ChQYs6BRnOhIbbyfJF0Go3dTTIqti++gTMfMm8U5/WybviAlzKQVU87oD0
SV1YCrucY00E9DQZ86/LM6R9uK7aZkQykYKcNrVgJu/Whj8Z0gzH6S951JtgnFkwjfEe/iojYD+u
v6CTgJGoiqNfwRSLlBQAVW56ZV6c/OJm5/qkTBNiT3O6TVayMLVhxhIlLZWkgezWXQS3TTFkzvcr
i4v4kGLgxUO+nsM9Yey7GgEC6nPn/6eWLWxNAfJkQoiTMnlQkAY3r6cWxGSA1yneBFg4JvzJ1CtL
N25QeMlEgTu0CigULm6ebCn6Pktqx2c+/xArao+R91rERMl0cvCeSrl9tkRAaF/soT/Triq+Yrsb
n8KoCoGi+7YZJMHzEEZjjpnxGnb5cE0jkyo6LBm7BTIr9PSBUX5sx5gMKVTL7k2dPjy9+FMXJC8b
rKWX4ZyydCm7OW1x/p0TcQLbMlhhBPXMzt8F4oJRA4pGfPCw3U7LU9B6V0h78zsVpudArDb0q4pN
Uvnm2jZgHseUbspq1ZScZAU5Sx6vO1xmyclGjMtuyrt73u+UdJipkrjVffkrBCPUk3HrmjOoj8c9
pQdprKjUpsQ7ufAAZYh3B/4cBvpAGX+cDURlk1OF08T9m65qyFi7ax0xkvg+0SzmBJvRkbuBF3nh
nqguhRIKnLbQtYteBTfOPcD2s0i6dJcR9vROeuPGDcXAnDkl+/nyKNVMKsvNqHDWKU+hklGdpRay
9tbtc7XtBhVK4IsKdkFjrUWHvy7CiXt9eBndPSJ8xsrJ8vvz0BqagRftjgAgtZP+03wXbm+M8eB1
TApUSRw5Xv3sCHV2y0L9+lboVPkITM8UbmRpHF8CnmUwz1C0mM9QN/ILDnjvd4A08Yt+cSV2ifYc
2VsufPiML2vdj1Qe2+61lnOrJeHYY9Tk+JbP8LqnrHaQ7SYGEc61/8IaESm5vVBnHya3RfFppZfc
C5lvNVdso/n3F5+rx1Y6WNQpTu3z7RX8erdkDow89suEgNZIe0FHmVPfeYpX3HZDTF7h2qKyw/+Y
b3RvxwC5V5Npj53EI47pjCvdgBi1hcGf+/y8vsTtbjhqG18lLVBMOalyb1rR9R00tv5INPuI5Pef
PWx8rnUVxht4MEdp2GLDqxX5cmvJcwMaZfVRoy+PXeRT/FJj0ATp+p2p7HMUMYVVvWturBNWoFOt
HG/fTCRCbmtrct7HUvBYb/+JWzVyCSUUEF0QhuLl/OlpJE3XpLLWjNSOT3uHcdv+k7tBeky/uyuy
y3L/y/ufzG0jt+XyIpYEohjAnMfIZpq/UV1WsRRipTr2XIYssOJH0oJ575YS0wlsrRbBJ01ITCv8
bjTZLacFG1Ttgzuj0fcX7vguip3ot4MsH4hTCY9IZYQJ5D/CqlbbTACzhKvNSGlCm/9twsWCHXQk
c99bpnSZ7bMyDtPIYy/zitbn0vGTY1PWCpy+f6Z1LHKUw7t14qudAA+PdsMKyfK8lb6mjAgPt16m
V7H2f/cbZH72rtQMzNTT4FyXEm64Haf3vStkHCshsjVo0r+y6ZqZLhaegjuT3MMsvguzgaiWRK62
Nr4JmjPYwMMSiJ0xRlyfFE2HLbYgVPd+xdmGAhEnqkBQogxdEhUCxqEB5qUp/FLNQjrRF0T8fE5P
vB47jhZikVObAs/nDHNc/ri/hZZlVvGCvv40Brn/WQRD11j0qkjYPhbxfbKQQ6WGLCYg3ZZaf9Fu
z8vkYFNLGwPTDJT9AV41kBHQ1Tc8vC/jRvcaYY44nJ7HBD4f7O3FYkIZkK9EIcyateLG4hx3in4s
+QUuOdMS15WdQctw6mKFAPGYSWHt6jpGnyKkNB8xlro+vWs6E1hriwl7KxBotxlb4b1c2HmEGM8R
X5g21ZvOua/4fyurxzff+1ODkNeCXT9+260hEpSjS5p04zeE6s7kk5azrKZA/avQDni0qbUrCUqf
wsSNzy1AASmznTaK9vt+RzJEERKMXrfmbaWoNYaikAgVZhC6NtKBbiIT8/koOhZGBXm40Vb6qhlP
faBG72E76WCXzllmo2zxulPvM8jHlLJjvZN12eKjyPYUP3tzb3znbFkclk8zoI/yKJNmkhi7qSIh
/qVGo2Q+FIO9H7yXnKc55wolIht6ctdltyybjriRjBlzBCL1vbSixdAb4yTDiX3ikSMtQO7LBkPt
vX/f7015PC9gElyZS3GFn7S99tWGlTUX203cVooFtoRcWXd01cuibohRECU7AejLT3oKTIuGbAK0
HuhQDIxgCOO1WLKV+468Pa/qOMQMWF/m50pz3LUK8gRJz+E3OW8cGbJPh9EVUd4/2h8Oz5ds+odu
AjLxCjEom482FoTOQ25sKUVWdePJIaER+mC7/nsThVEhY0MKd9iKythcY+K75iI90qlyFWC8T1kE
jyFhh9UiY7JuiM177EAusoES6nVeAJl8Cu7yal86piKblBDpnwgZDgz29YAQ0d33koFRrOT2HX6J
3r5wtFxpiBOF7DMM1pGAqTJ0YAbvhSJnFcCS10hw5txgK+6xBMA0qmuN9obV8O1k42/l10v75jrk
5vCfTY6mjWWpzowFGD5CXaspEtg67ByOPTebBJ9Q0b/tfB2T2TakyhAHQC5gkiLImdEvcICi+0O+
wkTVtgoI76WDYKQuirv/K5PUyNWro2YQGbN4RtyRA3jOdsrmKc91CfOAq8JulKAZde1R//KYLn2J
GoBVCewCIFWyPjEpmvf/7NYTMXxlPlCA9AiKRDb3+sEYHDUuosRfyMRQHad1Tl/FZrMhZVW3Wsk7
EmVwG15a3R0VqXK4FVvC/X10NhRnUkrsBN3zSVcgX13IvHWhbBTmxz5LAoNARp41PBvPkZUx4Caj
zVWwKE89A8w4H6SgKknIACMHt+AYBrybwSFVuSrqq9LS+kTV6jB0tFPmmPKigIay9q+GkWk43d6L
Eecxf4FXAWrbKYUwaLKSn3cRYS2RsLLvqpebaXc2hRTvPDgPlu5v8NCCFYVry1FATKJe0gRJSnWY
t3h8OD3sLlixKODKA3753X5TrG3la5TpycSXqC+WTaDc33+O1VUxnLMcXoJhH/WFD/0ya1otzKyM
qKQ8Vwngw+ESkM0GzpfdJlA9jQxuB13FDIiONaSn2fImN2lOupyv6SkY+UzJApUw5ebBa2t5XZgR
Gc984+t6F8RmrIo3U5eTyB9Lb7nPG9gOzyp6NIXIM2P3fbrZQMU42/9Kpxtf60PVp47voEzSc7fu
28CCg6YWA+9dzTk4ClnZqQ7aUY9N6c+EFiPWYyWckQPm2V4MknvA+ozmrFXMhSwfndsfv/cLbdem
+OaJCqtfdIqtuoPcV3BfeVhVg2tCXDMe0ZP8Qhzn+Ad70yZYTlROeQnzoEzmqFbCfGrSWzxtPHzj
5feQ3twWTb9v2IqCuHnfXhyuiDuOgGQ7knRhpOY1NHms/wdkLXVA9WuakVx6rc8GYYoEQi28mxqC
ZaD1B6zFXmn0poJrT7M15Cpww8Tq6aPCA5kP6xFUCoTmKJca4/oxUqY1FODl51DrvaNgENLoIcNb
aUyeFgnX4nxMTCKengD41+P1NvjpmIfv4D219dgAjKaUofZvwfrCwGO9dD8WTTSJN/8VeNoJN47+
PdyfTlIozffctGTV9lEXRCP6HC80ne1n5CwRyhnSMcIDAAjScND2tub/xuXWJlGWP+RowaVtrMJL
Stw2DuuIdKNZRZ1TZt+HoKdjZavJwfDxrqWIWGLzoUfK0KMqlu1gawFcLPtEccJMhlimeGG5+BdF
CiC9dEjk26AUnuYFTlvTSd9JRvYvPTJ/Oq1Q5+fJf5+APKCFK6hIW4nekPWApwI7w2E+QVlwW6HH
D56lqVEwattgqi69KDuJAzT///P96+pZrrnrhnQs/WZ/5o+UE862XNsjXyzH8j2nA8P2lZ4+rR/U
prH6icNV/+Hz1QHPXc9v/C26Kju+SQr7uZa6yt2vg2YV7FZ7W6wd7PslhZ0kqDQyKI3T03O8tWQN
PmbDYsDzCtOMxY0MGlVfbESTbmPmveAfxSMbADo4WKA2z7lZlQfdLbFqkGZ3X8x/BpVBXZjYl/hc
4fSpdWUsQivy0hEFni/7+AWWRICfXzxlQ3Ll4L5rqzBSDmrjn3mB+ePTEr/8SZORCd7yaLVjIrTx
LGb4QCu54Ks/rDjqff3rkZ8epdBZS+Xc+P4VRzC3705XRX+aeSJm4oD3DKcA4ddK/vJqQyOuVCAq
Dx9Oq9R449xa+3+aEDWGSIjpDH+Szz6NaK0dszVpnN9gD98ZaDYim59UMoG4nRzP1XP7dj8IL+ki
tik8fJGQNhGgzMYKGx6lx1uvnBPyT4JfXhB+/Q7dxLUvF/sRoqW62uFQrWNe/jDU4OwxWxciR0TZ
eT6OyjvzDf5JvEQ8xjQPO1smzOlriMir3GhvwJLX5frNrP7JqPHqAtmZPDlh2LFCtS4yMOPwVsgv
h45cOcR30eypt4r9+OWkkEdEZgjGA+b6883mseJctqFUA8CLPjQ95HD587Lhx8MhQdX3a35gsJoH
IBen6t44ZI/CFHrR1bsTxew2bpazVNathmxj+zcOU8E4xBLgtTg2d/ApBmninif131ULQMsC+4tG
+gANGCyB9sNkFEDL5/1DNROsxzcBFDrEAyzWVqlJvHmveRF+w57ZBcd97lgnnHLRMpJlJCvkcAe2
JBRk/3dMWXrhr2KpSnYw8PDczuiq3Yf7sbCgHrXZhEy/QpkPVIdarXUuDlZflVDXabdZXEEZvHPw
onM0J83nM35kTAY80G8aodF6lAaboJHcPzt1H0QZKwR9gd4VWUGUVJkSIeoIkU7Fv7DnrkthUhYS
Lw2QwtU4u+qJ+pLLWh9FVCTwCYUkUnGvn0PebRZ6HoXfW5jwY8UUj1zaBaYJFn8M0UZ9HwLCl3FR
A7r8G6tRnYYBca4hHisGstRsOeNarYDip6aF9+JrmOOcnaLMP/OdgQetELz/GWQpAjEZBDHC7j1J
DI2B+L0/sdlcVpI7T1zldkDZ89gYEVoe8ohInvT90yTO4VQPJzlcgNM+V3WerMAmZzLlpeir/eTO
6zO/JOa+pOrJXwr3JD00VX5dNo1j+1WO9yp8/xHNw2V0ppgaklfX5HobnkiZg3oSAex54rTMZdA5
i8Wu7z7e7D6bYMFt6VY7sOXfKv38XReID7k3pwCxMIuij9LTEx8taKeOJ9y6fSiqI7m8H0Q7Alv7
nCNwd/hCfjeFwG+eoBRh6ZRyIpbj3QcYlxK0g39b2aXOgPmLDFftrEq2YtogX3gUIPumNuVJyi23
wgsRSUKf8KKzyUE+kqgSrrXr0pdz53d4jGkP1KKODFKsGiuihxp43Xf5IjBoNb+9peOKObs0MITB
OcNLX2Ln9ylyWL9CnXjJono3XBYNVAhGEfQLS7JEauGDH8KBYRlAtxrrM98pSz7sGmV+F52Ucj7T
OMcEsFK6BgTXF58gRthZcF7vTAiZMRSol9rqQ4YHEsS0WgQYdMCyhV+t+NMdKfqLh9SMHWjgFLme
oOJwr2RX1L3qMrFrk1sVxmATv9DhEApimmkLWag7vxHpZlk/FOe4SwAflPRvZ/qFbGnPDL3dNqI1
BHrnOMI5JgxJKw9VMkcJj6sjPepSdmnpdUVAczD3jeIA+ogrts8rqZNn9cKjP3V9DoNCvl0tqHSn
QZVt8cwd9yeOYRdFrmZP0rkIZcP2OHko8p2BGY5S/LzsQZAF7XEeO8kT2EMWUQUVvmEG7jnLOZvY
biU1hM5Ufs3GZ9e2xvgVGI3TR6Y34Xfsj8Be17Vw+62zYJctg5Bd0V63lqtn/C+bf8Y6s/RL7QiK
wC6jRh78wiQKA3SDrg6XmNc71dPfZMwEqHRSmxZTsZyo7IJkMMh665zT88kHUjJHp0pGe422Ckho
I05hSDMUok5pyoch2Chh4FVHIPh+uyCOnMYx3urFF439waK8qzqGokO0hgNeq2yHx0pfMxwrjtUP
+U1cQbvM94KinD+82PNischIUYCWkGgbctd59Rr2tSQguj9PZGIyAk7rorcwluNEZz8cu4EX2tnw
bFBrhh/WkWWD4ePqavu5pAEUNNBngoxEo+6TJwaeUtxOIppUjAiVShDPg/3FDr703qCskbwqYDAj
9guINVAo5O6ZFLMEyOmIE23Kws5PGcFx9+iUpSf+2psmx0l9DM8XOeIVP9jvB2pWPDENKvOXjMLy
QmqgCWT7kjmvnebVcK0arAqrYjAwN0a0OX3W5V4BnYhyeRg6flcouOeUx+GcrY+ewuIWcaMcIsn/
E4ri2vmy7HYOgpjyTxn0l+bWIFBXTyrC18pbc16WfKQ4rQ+j1e395WrIi4Z41ZOlsowK+aLtcEfF
1Qdz3Rxex/4y0cDe3uZIgJh8G2pl4LTRkINpgYf781rk6u02/42axMa6Xkw6yx/RFbqQ5FzIxog0
UonTiGqRnLWY76eCQ3KUINswJRgJJH012RT8PLohCnI4P1K7TVG2zXoNeLLzWClSF29E9Jj9hkY+
IjffcrqZsS8fmZm8SuC6Wb5ERmMitazmyMco10GUaMCYDcVZyOZkI1/5/zLfki0gnP7wpoiBK7KX
wZEmIySkkYM7euB8qZh0YUQKluwYx/7yJQfJsIGnIurokuHwDNvsE8u0f1nMPL7OkL54DXakY731
HI5V7AFAmTM+e1cABYzd2jQSlDd8F6bnae/BvkQCf5qrKFBRgNb6Ra2sbZD+aQ115AXlAYqJsYKd
+tPXg5vpfIL/Hlk7DwjfCh1XjAy5PsNKl3MN3X8/BWpR4tBwdxB1tJXZaRgkUnQ/DuQkjxXAMBoi
ROj0YuRKsTv3V/q2jHqznkSL/h5IVtsRg2A7o0UwPpq9TRnYpdvlN8F7C05N3fqWpyOmAXLqh+ox
W9HU7nU8h8NODVUKbOX/KfMCa6a1p3ba+8HHtQcZ8ysJ9Srk89VACa+Nk2DSjcneIIKoDUHlqW2J
tsLyZp3immcrIm+qaL2gjp+aFkASZ022VfLfS2TozMT+s9g3egB0M8Umnzham3WT5BQq05Woilqz
DbiWlDPIZebz5/0FUNoJvJ7dEQkCg/C1nueU7xWsllElDhfMjYwt+L/74yqSlbpd+uM7N2swQjm2
xipod2ojB7jBciH7AzTIyV9yPIrk3mTTQ6JniQi03UBxqcR73J582jK9WRHvqJkHzbPoQjvJbM1w
k5LkfsHWOzET6dZyhkOUb7kDyDAmdmB1Eoe9vn8vnBO3RJV8gSjKgm77oEZa3sZL+Y4Hj0Q3ruYM
oukjoFQZZ16NGK7LtLwkPhSBli4Hy8P2CrZJ1gDamvSeIUsSV+ZkVRA5P4wgtmrc1V8EYy+nMili
wQgqmwzMrfiVZQdvs7VRdMriMlatwFrX6EzHinTKzE9Hw1uKrPvRCndsVGFjMey1n77SKUsybrwB
a9Rw9JNrPVGyvCj7QtPAaxvlx3X3vFPsrElLfiBFAE2udv/dEObuOck0KjRBiazQUIOZZvATNguQ
G5vY45+Eb3Um9eLUbshBkQJ408G/NOYZJcJwWjwXq+Y4rNmt7zI3TL42ITmt3VpYdiXO71M/YGdm
DyuIcL4N0w4i/vGZsxOus+YJDw1eZxf5T4+y7tHqRaSaiszfzZfBdLWrfch0SCotipUD6tSfcrlJ
tZVf1QWyVoSZk9W0oOmeS+X79CNlVDpmYt2vZ3C4sRuEcnioi+WzX9Hzfv4hsnThG7Mex4gaOzLQ
xYvvAUjamb86YmL0sqb9EkpXmPXJEXIUYUpoqPZIE8eptAs86WMVGfUypB+tJiuCrSIt2+E0xFt9
L4WUM/kEUZyaQFLmsQ2TXV9ZZ2qlVL9JaOXNGQ2fGY+6pzXYskDY9+31rVXFg8OVhKy0ErK+ghid
CH55RhmsUpaZwAZ2RhIGcMykel5tV07BJHnRN4bJrUoEwUqsyQETRpPFhSv80sIgnzFaQGr1OLx6
SDjCndLUxluaFd1r5fEJrYLnXNRrVKJ2LQD6qK6AIjdBk7S55wBa863PQnI1L1NgafdiyFUHoaY9
+MRzyYL0nUa7bYqJASc5UI3jk/xyA3P1I9Yi2Y05oEL4gLUN82zXgZt49vEH4ZqvMWPq4kXE3KsJ
BkU0YpjkbG4CGScRSqd/UiyFMYc1307ontBAzH7pFNKs4qNPMR+i4X/ILnRcJhOjjYCCkRhq0KjT
2sHjad/o+t5dU7pvElhxwdZRtYcqa2D0fEgdAaIXSr5DT7Cg/6HFFr1iqM7P1GaikXrlCYKPEXmm
5CQB/v0Q4JvgyFboZDV76eb/rX2Eu8eZFI/qZrkpvg2/6YiQyka7o4FGwxgFgVun0gvBPjrPAwcp
xxKDU3DbRvM5HqI8PjKNhlcfQ/KWuHgTdYwciZYDuGCpHeWrWGH5D7tJ/LXk5LLuT6WDNtLDymqo
k3oXc+1M68X1zzpSrXKn07jy4INkShIigtz9lnvVJn2dL5pyZdu5PIOU1oYHFQCOKlgp9lxv57Fm
VwxARDivlTv6zl7Pe3h53S5y4YkN9ZmytXuSlcpQjGesjZZsdSW6U+FNynQ8C2jovFa23ejjcWCs
hd6UxP9rQnx1E5kLDXUYarRrmYDdqNhXahMNKybHHRQJzqXT1eCoWAAG8akGMcJTbGiWiLA8htBJ
q06GFJ2zb2ROBO2peaK99Ez6YLe+Gj3aVl+zuvKvkNlQKmwqW0+ASWVtw4W7sZEn0avr/EXL8PTZ
XxdqkS/tVqRzHbwHkgPuwmT8PkQpUCG0+0m0QWq7piej7Hgesq3K/XYQrqwIo/Bc8GsQiAw709P1
uRYI/QrfZyHVdMfEeYAaOrLGWbBMKrFvAmOlKqczumA6xz5Azcd3LpuYAkaGCQOprW86dI7/n8Qc
A+cn7BIjwoMyU/xsrWYzVbXydyCcgUqsHRylAXOva8U9CrWpNW9abNFjnJUeqTX1PHlPRdCZ+GT7
6oI23qfggQgPZxe+Ponbh3BYsTRWSC9kZ6YSOhr28/vwDuKFtUDCKeib7+7Op+XFshq5UbooTA2q
Zo1tzH8bGtdKHnV8v+K8J5PisANMAFEYXYjaDlYVVmjsbe2KHMMxqF559b8S14NEj+WcURD+T1H+
vgESPrnfdfe0DgU8cQD8zp9aDY6CTkuy+eUSpEtXHKF992I7D+vmr01/bq5WmBOdklf5RPW0375L
mbneO3iSo8JgITUzc4STsQkcScO4fP5gMc7rXd77w9trvsW0lIexzOg44Whfqk3mv2C5TKxdYCSy
RJdO49X/QUVax1kyIYH8URWxi5I155X3bfseggLkZsG9d00EpiYkrcSmdgvIZ32aWvxG17velDcH
ORaTcX9L/Z/GgYAoS7Bpdcn5qH2CJU09takjOh+fKjXA1PSfNvRta4NwuN/6hdTVLrRFtQfDaGPy
S8/Eg9pSPI3cWZso4VZKmzdFwmz6zHlfx5SIW7HFOASH/9BPBdX8nad9rieg05GbBsk2WTxnqoiK
HQ8wGa8i7Ho1QEKb49ENEJeXlP/B2S1RB94ph8RGXIvSg+l+g0QnIPzk+9kKUfiBqK2v8XYNYyY1
eM/6zFVkFazWMIHCnLs0cjlaxLxN1OErtRrdOxjy+BP7LdOYqBnxNFIgZogw5UYiAY9uZ9A9d/XY
+PBHCfEgKkRPMX2ahYj2Bv/StZXpt4M4gXJDmV3imiFmteYXUkdr3zEqfaODt742otXXj3XkcaoV
+pkxs4jTUfaXXWa+Utsmn0TZuZdZlP5MmCMY32Qtm3cQYLFsI5klQO9LudkG+vMsIxd2mb8mVBoI
tjVwCR6RsXERxhH9xuZEoK40UUZ7mUUTtTLrooKq/N+6c7eUTN/3ETHlnaWosYg+0UMLqQFYKd5V
P17jr78SXwxjA6DLViG5KazmSgYjUkSlQZv2/jCH7i5OPtxrxfAnUyro95U1hPQZWjn4iJ2j1SjL
V/wQeA0NrIBQFCMmBSD/NPkthfXIf8YK7DSpx16KIBmAgRF9d9Rg8uELvzwNOhd9FwQMBa7CqPz5
NiYj+c7c8YcI1VDcF0l9jRXLxdzC1wla8vGIvrlJKAXbVnik+QM9mReyFENFYE8ondbvjRhvHv5I
RSTfuHnRFg6qPJd2hdchZex6xvtTOsD9RXOxfCAaK3Z9up+pyVv6tbJPJ6kOQnFCcuQPWTSn1Jx+
yMZsL3KoHnEiWegk9NJQeXsTlRMTUm2Hh3LV2GVG1mKBcTd/rxEa7ylmpjkt88r2wMSNbxXGVN9W
6sQN2jGw7+vvFsV+1X9P38g1ocwLKfJFCx675z8itP0tMLzc6shAuWCkfFAoHcbY6jQEbNTvbqg1
FE32Pyjz3GDGeA+zDiP1SpT1nUP8HQ//XxpjN9ul0gQZdoag5KTgtf8K5OLT1QWevZ+1ZyxJ1wEC
ZcKwvTmcL8hAl8SeWnSbO/1ybcqAmGy5Bxx3cgN3vel4MttKA7x6GtvizLfu0K7RyPq6cD+3Gepj
r3sp0oddFnt0eTogF0dJ3hNIeoImBQKQX+bpWcDpCeCxecx8qhjfcuuYhmcz0a+eIKORwiSY9Y+L
QuVDSLs1tgKmx8rXX0bqXT1t9HV2NhhShy+nzYp6uVseuU1tqWQvDgI9Ar7CeI0DZX3iE/ArAEtY
ClimJQn8X1AIeh1ByLQ0fRBZqzdgsa4zEevn99p98izdKt2B5xgMkg0B2V+nPVyWIWTtz8AT53VA
w0UU4Yzs3MVl10tKhjWYOFlQk0x90262dO5AjUJfW4IrMOdG2uf3vHABHCOS/gL+09kU9plRlqhB
mcUE92CaPAaJFzs5jsZMumZKu1gMoYUgc8Q9r/eSEPe8rFFYE/8QVQatfosbcFQKsITW3mSfoEmV
fhFaSGHyhk4Q3tT22PJjDRNFWL6t75j92+Qp5n+cP+SvcGxzWeV5Vt2MUd/VdmeSDbF1JkJLfYnd
ExqtmVK4ArUtgHONcroF9pSn0jVRuM6EQBproutJBHBje1miFuEZkW00jD3ghZgOfw53xIS41Grz
y/7t+CZKuy00ezJZhqnP+AI31Xpik4/9PQHtsQCZeIu0deQ7qaEIg7Zr6LBdmg8QP8ei0k6pS0Vl
4iregAf+T7sRKF20/JkFyyM+I9+9kJJC2qfdiWz7ha2cgP9bGxMFLfN2fsOlhbrnu+I7ah+6qjAv
MvqLsf9d7jlOV8zsO79an3Ihrp897oIJmNVQSd57vb8VI4gGrwowTNA+1cxwCYlirKVaWauz8IU/
6MAClVw1L92MLX/uS2Dzi3VdwSImk+2Y2rH8LxUM4FixR/4d+rALKrgyPGVS+cG9zTZgMSYisphK
Q/XolzZQy/FU8coNNaYCv6kcH/hQ7klDrcv6hHar/ebCzplxGHMlo33XImhDRNirKVDmxuTWerpm
ZzaGRg3ldDjmA9gBr5yz2bU2u79OaneNBc3/lB4imJOe2NFVvqT2Bq39WiVdjlyCgTcFfAy6dw53
Y4YlMaeRgVTijNwGzuWx3Hl21Vrr829oOhljkM53+s3ZLz9qtY6VewyC0ffQMkaW/E95pUBi7Wkm
dZKhP4XEFOFq1JvWZ5W1xNFHvLmO3DncBwk7vDlBIsGqdkHCkASySYZth4lHnFwUk+4zaCk1if7U
CRLBTSWffsyJ7Ylyfd5kDYeyL74BuJvWAJKmzPBb7fJkw73Yz94bW+1EW2KiqJHb6pTTRTyaM8pC
QXa71T9Usc+ABV1dZnCo7dYwHNFoBLQu8mC2eyGf6FJ8vrNyDnVqTZb60I1plGlzvxkBgcBtj975
CrhqelqNsjq3+Pka1+LZQLOWV8VS5VvTTWLMhZA2ioi5D9hpC3GrHa5wDl3U3MDt3D1FQNCGq8a6
uzvzi+wkXimdZid47gKz398BZ8XWQP/+nBwpAIRFzzb6CGtek7/zk+xXLCwMXIULseD1X/Bm8vVX
4Ant8IrG61y65uwhJsH9xSXv3h9goOLiLNag62BiHGyn0wghMMDlU2/y7swRekrV87YwkE1f2RZF
qhqtPlNCi4YMW5+6Q6iFHRNgm6wSGGU3nbFtO0IQ6J7L0u/TRM08a9oBPvs01lqJjrBPPDNSBboK
NH/Sz+1H+pb5iH3r4f4ryNSphdZESSj7Ky0e7S+GZxDkz0FA/Cu+wvrSrUtUi5b5F2LBFhrFgvSq
E5PMrw1zJSlzwg8mk8rnu2DpJVc605xgu+M7zmiWAHQfrpveXx77vHk8E5PauiPYQ9BYtUdXFrdf
arAaNpDnhuZtmCHYZLQR/o38fQ/qrV7EEoM64Y8B2SFExySzyQ40OXRUYBiW1b+qLmrq5mChjhvJ
iCqoUf496mxAUq0s7WzBSjGHnbhN3yF+u4dGqI47+0JpNo+GFyTcLcb0xGCyX0Lr7WVJW9DTUkS0
cPXMczf9KuYGCom+gYn11vRfDcy/5VOOYy7ZTdzOQSeDeRrtrk1vgVt+1RBxGVG7eyaljLUwQ+ye
xejeX7+wC5AL90EJS+E4mZ2BNQLWqQ2h+9Sh7bFAmlntgqoVXRLvM5x+5a1FXjv24Hm+NCyc31gd
5Sk4Xxpv90VlggQnwEwhKMdzmkTXELoQfw25DWDaNuEDtyJdZk+mXF7wqCwcEIV5tGabokpLgZW2
TrJfLTkJ7ZH8tEeEHCGMIOVK9pToF+zn1slpZ5Vj671WrhQb9Bw/zKCX5liET3wIM1aoL1AX3a1w
ULrDGo/WW7Go3BHUp9/NFagsfyZ9Zt37U2dbmVevYLJN6W9F+37K4RQc9hbExHO7JF5gIaVfT/Wb
DSqgLylHTUPjUWkKKDf+QCv4QH91zo7Yc2QLWdxe5i7fFbNtviCsl8wqf+TF/zyEZ5b6pPvbTCu/
oNf5CVfX2eoqUuPmjkUptNScetK21HSLbTkx8T3VQvE8llX8L+/hj66G8DTFpf+MeP+V44enAoM1
+a9I8gnmdma2Y/eOxohy3lR93cYeX2pYF2w+piH1R5TNGsJr2ephkOCO3F+qrKKL0kGAkIGPRcNK
MfOerqNyn4bRvVUreHAxpgXfJ3db1d1VjBnXzk23dQQ+MreuSnrPsWThFs2VddIvUFziNFksexnV
qKFuVrGTAeGJUllayH+uxlho0I3fkYOCA75BDCl1Gw8hlVirBn0XbUDdgf70o0JLz5CAKRV6W1EF
aChxywy0cXlJlrPCoY5n0CBqer296DKfjrM1DIaCrktji5oOfOs/kGhP16uq73QGuq5md38o+Kpz
fFZwHf8d5AyTr3gIHbluAfZYtm5OC/Z7v7xdmEoJkUBncETb7DBOlXWOJGmbill9pCTtRraQuNs+
oxnR0ku+6Z0Hfv2fli2KhkHK8Rw/ls3gQ5DPKmp2mdumFDsqn5pW4rmdUDVJZNGAkLljCT+QOTr6
We1P3KknFbuJrtxno7lDMwzk5PI+R3Ddu0UjKnrwmuJgzB0TmsZeMqZRNGpGCzAm7CgbvYIEu7r0
4HwXUn3wISiINxpGDs/JxYx91NwWnlzjFeIBAQvQgtvSQzPQfScxnT7UQ3kERnk/dwqNKfOjvpLI
Ej3WB0R39YhtCSlOZ+PJl706dwx/+NlL7IRvYHLUhNPE/7A5v0t7vFh0KBOCZ+Mo3F1X+rJ33Woy
BnEE9cCGLA7jsF1P56mtmvthqHrGuH2tFARuGWaFb1Wy8MB7Rsd1xEdEN8RDRtbEsULm4j76g8+M
HnWqvQkBWvzQBTYurak85jbdZ1LnJ4GVpCyNMDUozEKIezJPyKziKPkrKNXMv/YRvs/pAwwmgbv2
C/VgyyU3fdd/HEKiWQWqlSFLbZRixHxZz3gDXVWk+vwf87LzqH46MxnrxNpGvSIHHwh4yxinCbFs
VUjHd+UaSYsxeyrU6azcln89npkpox+DXv12egYMEiBn1Va9pfY6cKPSVMA8phLgeECJPnDlPzFn
MjsgYbreEyD5NNXba/fa4+I43+pzYSrLzio8jjB9vDP4QbJ9eMnK5a60ZdrQ4oirKRmOhENP8Ib4
6L/ic63jjuZvaMD2ORD/Fsyfg8RHUtS72waBOQXCBsHwjAyIC/hbgzdgnqKxUMNkcZ5cn96hu2lZ
x4GLhnZmZy52AZNnUSIGY1zJwUb1XfWbb8ykg59G5tJUkpXo+o9fWCzkfZ5cSc67ccRNu9twyO9T
+wyhKo8e7+KwQ55S/uXfucDqVCtcl0VEFd4JLvnJUwhrqHOESajcTz3qoZgmZ8uR/e21AM5Rt8jx
FFPG/hInzcy8w3y8gb9RxSy2K3Ft9yA9cnd0rrdOooD1CQntQzbzjffrJdPfkI0BEh/KTXdX71hq
0SKK83wDaNUVCi+XuZ4FBuN34fXfZagwOQVnAXJYG2AaDG6wzibaPX3INrgBWJFqcFtDjKh4BLFW
dKyjS6+NAzHexxjpBj5Opb43XYPSLIEtm39JuJC7ShbzunG/eC9KLa+it76+PvgeoaxVtCE47Geg
2PfQ4C6igjhHvydg2b+UU8XI5P2/4esaJO/DXmYCHACbByaNFu/Z3fSEWzoBaOVSGHz77Ct8wE0G
Qv/E8bd6qZbju8+Qv/IIFvTeeQ/zg9lgd4Haac1FN86YcAbRNiag2S9kPM/uCKvgtSZXH//2TDGk
8gj4awd6Uyf9KH/exCEFHOka55BBqj/lYTq2gYkxqumDUUElbME2BnL97SHbbU6U9VTtO1VX59c4
XKFpBkMm9cAz2Z3MgWosSma0gGq04EDt99Ed3GmYvxN+GLWdEt4n8PnK6zXzh7Lq7W7e+ezkpbYg
KZyQPY8u0bZhsVDO9LPDaL9PUUrQpwb3RbVmw311zKj0ZnphiCYhuipzP9gQaB2L3pctH4jhEk1C
vyUzLw4jEEn2kAfCv3krkuTxu/mikCgTbhJCZvdML13/pM/0PqdWqpoD+9WdX59dNkyLG5bqwPPg
VgQr50lXJEJi3FMgBhw70Izy38tmXj4eQDMMElv0vn5tw748IebC3L3K1KHus8zdmes/BTpGyGks
tsx266mpk8Co5uhbvCNkuW+GPmEc5uVkbvKAliHMIuH01LZcp5DTo77AyrxUda0WZ4cJASZPJ3gs
TcqU8V4al9GHLHPnnTyIted9IaobYHeMyYm2JH60BbW/7XJjAWfR0ha7U5BQ1XKHZwZMQJOPHHdA
MwENjNo/UKpgHijRFNBQnw/hIC0NQn2DAKwVJWzmIW52MWHvHaxTmaV3Co6j509vdYDUJeSGeWdZ
UtqYezf7VnPqUGBUYkIeXrrnt3EWvJkBceuhbsMyso1qrll/ly6rQ/sKVEvlG5KB1fA6cBH5DXxc
2nPzv+aF3vtdAef7Wce3fHj+C+fTkuoUegVY8REb9uqR1LNn6W0qVeg4DjXuI87YVXKaxVrSnEi5
uScIZw0kK0R/SNtEAEjqMBjqp16RYasHtsFqDqeEL0r1bserhFJ1Oy6TpTI/ge9xQbyfGDn1PfCX
fX376NSbzuo4UzWixn896p913Uh3iJO5FkZ9yQWe77G3OYdmPsd4HxCEK3GW7pTsIB1Bo/1mFe/k
/X9LuI7pA5uTH/03+hpoJvvXmwB6iGjWgN04hDU+BEw6hfqvi/VWE1WJ0MAEy3VcbQhCAnNvpdK+
JntU4BSU/f3F3fysA9wPCaP4rNHsuRP5Oj2GlaXCM3sfN3+/B1qWD3Ia7n78LByqA/0Re6Gvto2q
gzVwJR3TiHciH7bou5YUBrvBI7+mPeDtcS8AUqSoGpfkvPAUEKO13uzykXWt+3ql8CRtI4DGSLny
bv3aDFL/oBJ+XA+JS0qEXR9uhWQ5lf+yMe4rGzs6JkN2T359hGN/vXwniyx2DJmF2UgcUnwlUQjP
FLVAZGz5d5Er2P7Iu79MwLwIxWdme294r7NFnQF4iqgdrKGT8KYLdi3xruq+iSqh1v/WNPUVXepg
hKbVvjaK4Dl8NUymnALKcXUBrvqLiQo55v11+tsntulSxzG2hhioCwqxjoFqTeK1W/1ocTgn+Jkk
vY6RparXC6yP8B8tNhBejvcrSy3vEvhQaPUFR+S5EULVtasczecVDjHi52PkWoJ6aWjHTMV3hrPb
AvoOiXao4Ud1QbmCfikI+74SbHoRf7nroTPsA0x6RA8YeSqXSsuJfCQBulgYNfuYvGOyv4p9+Q1J
iUswjsCgwwQfxWo9GLZzLG6czaS5tDuAR8KAvW+h4SrLbSt3bQigQOGUU6m50lPr0pkMducej/Si
qumny74VXlSJo88HSHOp1LKfGQ1v2d/O2G/WGuC4bQjgDWt7dBJ/5a6um65O3o3d3ZHNp57+wkbx
GYFhtnS2ieot71hsIlgoNdZVKU41sInaXbRZTIkSLVQVx1T5A+1IOasagYHUUFEwXLRy/sSCHPxM
cjld/LA6imwPvLiZTUa+pvLPg9TLh8yrU+vAnOtsnqcv/XrXeRRq6jcL6rSIMumVjJz21uk3PvWT
kemC6Mo4kqq/vQgfWnD30j7AolPGe5tzhtYJz1sy24h3H7s8mi7CRjBu937wc616pCwxN+BIsyqD
RJ7LHDQdOpzOjntYUeNzx50zeezuALa3LG1RQpQsWJwhu6z9sTco6DmWAW8MHObbTOyx8D8DqYGB
gByOS/TfZPNdX2oVGoMILJYmgmx9s1MjwZ5hGLSJLXWj1NRsGD+uh3EqG+QDwKQuE65BH+5Rq3KF
olr04+2UxApswA7eTTsBdVxCO803oIGt79ALom4VTsLrE4PMV1lImtdZEnZMDBzaGunZUG0XQgzw
ga5cFUEUsrz3vlPXXl09I1+JUghqR5UqnZbHNEOZmRO2ZlRIAy3SraxWrMObSlZP+L1pf29Srx2i
zxMWrdJLU7MmMqHXCNSWL/rZz/4lzmsx/CkbFNtwvfSoP2jnbpWcfp6eoPVSsiI0BihZL9QIxlWK
JZbI1L25Jfo6SJR0I3VDGnGk+cFPUwKGs10cYVt3bj0dnLmqrfNguB3UR4h+z9mO7LtE5ETSPTCE
+DmabWl3LIBEJTxq+cUQso9bux/Bt4mKdY0AiE4U8XK+K60owFXeTTmvMQKh3WTID49QisEfZ1E4
GIYAmqKfrLDmmcP+b6MDVeuPTI4WgnAIBIp8moQ7oIeVSw5h1WW9bY3GJYOGYtsfF/SQ9r3WFlcQ
3eMGq1KKeEIvY/s2cEqxvmwPLEG97UMX66QQhvEJrCM9n3mD4IGrxQU6hvTZk0ZrJWg0MmoqbzP2
2GmqGpvfPSeRKhQ8EnuzRdVN5iT603vdtaIpkve7RLlZNnJSuooVlA2b10x1ySD3by3gvvtfX5NX
HoBbRjolznYNBQUrOvnVLfddiuuac1HpIan9NDdhGLnFqeta56q9cTZOBJwYSLb/leidDSlLonog
BV6hfQkARmaPsh1n0Hq2pBfXSPYdPLRy+GxXhK0agq+C+TDtp3LLPRwKSQhaVdqAg0hEjXGAGgh7
luj0OxNA0bmH1+LHFhCDsk8fJSydKCnzwnOlMx+Nm3j9BA6mWgQNVcUPSojG31glMkok7PtmBjaX
sRBV7aTeRRV9sQ2DeZGQj1Oicq6gxldXirDxTNyTpp3Z5Di1CeHhNS4/lE/Chn9Sr+C57AZBuui3
Sta4m8PAQ1sthLA7USq7rjNYHkU/y4PWFC+rivAZSCLpjx6GAqTMLm/fhMUrn+nFC+gHx0fX/9NA
d+V9qxHSXmnF3ANkq549bkadICGBEOuRFf3RWnZ+uwGmUZwSZZPTDcr5T7ssBYsh6s2WQwqElAmP
r7vighs38EPmmGX1qzQBrVCQ8YgYGtLVJNr/0k34zT0ePj7jzNWpEBbB6WRdcdpVz4nRHzbRYWiQ
pM8UdTEPpLWkLCo8eUrj1Wy1AoiwTKI578SeEa0X/nYZBgKCHb5QkyqJVobEwpOOQ3iTZhpddF0l
K5hLHjxDqYrePVNBjoc3hqXeNjZL3SaEJlmgVvnSjjJUTgn6Rim9ue5eRQ7jIKNtdasqX60NFjJc
rxCph28/jot11gTBaxWw/bLjiFckrdq/os+kA8jI0Rxk7sxu+coL4MKCCagCisNwXT9gz/rGkZPG
YT5jb2HFTaPCQ7nM85Wy8j2On3FU1Qc+oBAJoFEtlgRur3p9QY+UAPe4rTA1yOSUOn5XS92p1ZT+
lI7+LV7pVQ5b4u8PI4erP1PVIzrCd/TUqE7s8wvcDSrtK1nVEFfRYfSgnnJEMhelKgarVKmeVI3i
CMoK75hmKqn4hTDODc6hmyC5kGhKVSz7/R7z6GSoJWQfJUzEkGYh8bGkEW3iHb+COj63B/LLzREU
CLb8ZKUBVH6CoDEqy+XLqhue2fNR+L36Ppo+Kc+ZyxNmwuk/mJIJ/X7zYbB3xqRehzDq09+m7WzV
2AOtmqUHrqNVhngpkW1b/AP5HBAqUapUaIeJPTaMj07SlclUVfLdxi9b8MeOaFN26Sv13Xx7NYzL
ZsMXIggD7RliaCX3erb1Ncjp56p3JKfqH/tzKCKOdcDpr88n0o1PHnPDVH3OVml7GoYktZONqir0
7IAhA+XsFjP+2/zcqedTS6YVoe/WfqR7C55kCHqeepsYIdEfkRxaVNIVIYvGK66sxX5E9oWO0L5l
chdGmNR6lw6PtmjG9J0EKG4yBCIaIECK50FXxEe01q2E5C59bakpHwC0Mz+3wkASJMAb8PdplX8d
2B77+CfUNgTboMcQrYdpa289lc6X1Sw3HXAiGlIqioeP7fdvCE/Damab0Du9RqmYtYXdJ64eqyZ6
oxBJH2wRPDq1lYImhjVOU+shSyPYosEdaMgPuwNk1ejeFtTRGTF8onKv+ZE+/0VYA8umWlp293Vj
zaX7OttehELp0ZXBTmYxdxr3ArjjN8eiYAgL/fWI6XNLKZ3u034G6lLOnl2TDtnP7qn6LnUFXdf4
fGRf8Th5EhP7mdYvjTaLVvhhZtHmbIujcwzgjS2eXl/OugKP4mHWSOXVh06fVis0GHXh5LFIH+Wi
sbQ8Vmf8vy6/c34QGi12SLN7pKKKr81GYPozyqKXEoC2rz41veZuOLH7z55n23eNfqcjSDyQjar7
tyZQcQ5Y9UrennS2y8O43BzDWWeGIAmxgB53KTAnz2l7xW22mDvhZVvYt1331z3axmLlAxniuSWd
Fod6n9+tJ28gBvAhmSta5A10J7aHCdXpmigNd/MaZspyMKOf56inuRPSvx/YGHaLYt8TT8xZFCJ6
6+DHzY2BhbMOV3XHWESlGBmFbgQdclqj1bz3HuP011Fi6/HPEZSGtjfix8q/UVOGFrZBUgwyRSJb
dYjhOGseaULnDOCL89nfKJBRPFytLByROwERYmcxsuitftR2zMcNoK0i7WP+FaevFT9gp6XYMu5m
pjk1jRwPu7c0+/cnzRnw38+kK3BZhmsTJp4eB8nWehedFV++moNKMb5q0O8t0fDZ6VQaM55x6a2B
2L7o4BDslsueVTwUR00QsKIYs0lAbSbKFFbYp9vsrtMs8r3EuKH26EgX7JIgBhSmTB1j1/5uBVWB
gVIJEjeCbPUnFeFTjM4j5jtxAFKwcJKQmVDujdiPlGcLP8PJKWlOaE9cqpG8M3lbugbhBgkNy9MX
28YDWDNSo5lGMasDl11lPinCWjXXRcEmUu2LzIMKUugr6G/nZ2DtL5/DyXRUuv62UhHcQEwqJ+Q5
X81z7sDdPh0oyEX5b6X6uajBBKJjDUZa+JisHNwScYO0/504BzA3peI9uowMw9HK9TjzjNOfJEaM
N9miVfJEH43eh6SdoAAAuwX4aY0y7VeECh+VNsFlMw0M3Gob2mKQHStWUDw2N+yDSaejqFhzNr7A
wK6RE3drXM0uxSsg09dAOPZ62QY2JnZ6zUpd5PrfvhY3dGU0t3bFTVSdPpWC2cpNY5fFJ8oLyJtB
rotHF58Oh8sqj4v6U33uAD7HG6SqtkptbuWEngee8uuFBYHrDbKGC7T263wyz7clLj0wwdQpheAQ
eU5xjLK4qbD7RTs/1TBVB0pBDArykBousCw0p7QjBhlfnvTLTtOrzdlpLwuqtlZz51lWI64qx8z9
sd7Ck95rvYGA5VRF4eQBdVnoxcC0eIPu22x6sDk9hZ68OdBzuObaKlADdVw2DMtEJmYJ6HxCsQIZ
S+QmORgd4PpqA+i7QprJiN+evOwOYdLmms3lAUsdVyIDD6FsSIWG7f5UXDwvNKFwcTmlgswsHJnE
XvnmM641J/FOFcNT/GTF5a0lygywGQ4aOv7+rAyKrXA8ccbBKm9VJOGj3Wxr5O+FjwPd2UMft2wQ
E97gGAV2mxR2AqFk9qWpNx+7qIStAsoGehi6Ymqd1idYNy5j6AS6itsSKSwXdRCY4MHNvGmAEgq7
ESZcRo6Eo2i/KZNy8kkyovvcEiaGuUUWCQn25lXQZHhz706ROpXomT53FnJKeO+/LVjDwmZWbhwm
lzTecLPYIwtSRM99y3TaUMqcSHTTDrvHYHHmv8H7x+YzpMWfQQyE0UIKSIP+37in9yJoDNFbs/MX
MfB+j9t5NGLpBfYicmIoy2r9dVOZhu0c5QebTGhxiyPDcobUCykNbZsZ5CMBymPD1DxG/tqJstYw
wdtPFBUPEcE8B4qiD0beeSp0CmC8FUJ2tBzx+E0Q6gGNmH76YkWw5XLjA+84R7L/4/5yAcl9YF9w
znHlf5xupnw2/lX4hKrkHWG9QnKuxYDaJGWh4OjeEYM5LNisorKmg/XgU5C6JMOvx9D13F3tlZ1s
1wIAtJr6gdxNZ2LxMrbkgzLqj0u7Aud7mXfDsj0bVdggZ7Jm9V/4v1J14pDa5Uv9gRlGcd8Fnc8z
VMHRnRNJw7jEnzfoXDbdmRCPqwCpQHr4UTqLU77j8AbYR6jczItUqukXsgYB66D8RGrvOSwGwCSI
wso7XhVZEQ6lZnMgZuGMml8xiB/RJ00G1nRcVajnZ9FF7g5iokNQQ0nQXo0T9ck/eUWavavCziDJ
+lrdxW/2v4jxHN/Dzr389FJRos+JcpQCSoBKnhVWgMjF9Huw4AX1AvzOSxqW5BhiF6l/AZ91zdpb
lDF8dVMNvF/LJFY7TmV9zZoxo1b6SfgrqUO5/W268GXfgjLOvNfVyX+6rnH4wZsvp5DxYq0atblf
c5a7xqXL162ABRbpOgb+IuBOCExrWxkaJ2WxHdZL/zzU/CxLHuFsegzImD5O9Cm8pEJGZPaFwGeQ
dbWCJeDU5yLlQchd64kIlny0xCg5wsqz0au48l1sl3YBqNFhqE5Vbu0udm0binOyTdzsDNognRQ9
3Qz2xAjTTxXRAmMf60jMYLyCSF3OOus5mn5uwv9pRrMkvICalSbDKrjoHo54DEatKlCJ202bdOgH
3hFI5oPu/2kXr424Xi6McxxLPKmbAvB1R13TFu4Tiij+yJPPA7n8bj1JVAG9OX73rizhM4ZNUJns
FByPGCELo3mIW/NxpepIJ+ClKOtSi44dt04lO/hpA/Vzp6Ya8faTOnK4PzG0jMOj4+IJJO8gyW5f
6A44ck8Iwop5BZhnwRAPTHHLDDVcQRXrYtc3uK+IzyQP5NQE5tLTeO3VSTXBOxYmelmlo4Dq+4hJ
zmFH7CzNUeUiw4NfnKyVQTpDzPHJG4CA+9OUBJKUiwRrvMEZORVs6ucCZPH+SYZLh2QwYo72QM4A
4KItJ+BPt9q8NTGlun0/G8X7K0sH9i3qU5UZ9gQTefzq1su/lvD7SGcgz+q96BFNsAXuGaQlZ9b6
SzmSWfksEIkrHv+vOw3lEYe4PfxPx/94jRuNg4U6/iejSH5iU5FAAvchv84J0/s2VUeIvGUs1zlp
P8fAApbifGcW9ZYrF61jm+U/Lf0fC9CBxaKpn2QbQGgNqto3/qL4KCND3hyZp/kf7lAIaZEqlnwu
SfXVblRcmxLWtVSF3YSuCo8Anwj6WDNP+3JT/g2rOuHDZluY+HLu+fKzS/mF8keSdnuGeNEglT39
8NVJojZiny+oYmFr2KuEpu3HxxVWsELcaYFTEGbrNQzfcWhFB6R1Ff+h8Z4fUDqxyIbUy5iohklW
A0YfUiRAspABkzQ1EDMiZMU+gaj+XQ1r3lfNbkJeHzwGtg4WMzqkwKpz+QkgVFyjwQZqGmjSZrRB
JUJUMzaneybpsqBQh9Clb2U95UExYSWsk/L1Tgzs14OWzGIYenbN1veFqF2VpC/ZJb1G0qWoCs+V
QWdNg2rN84oWKxNgizPjHJIzrfWe6gk8s5k20iF3m5wFycT5Fm2ITkZztn6ml7ky8JKUGOe7y9eH
kDS18xAwON9xbwoYc6GT0H8dGr6GOPk/DscrP6P557RXar1qJmO6AuB65nB8WV2fx8fETuTg2eox
t3a01YBUu2umbyUalrcyrmCU4vsNOSpp9tSWPQoeE3eNEjnjV7BFvoH1utVUsS1Qzx/e8hJFmi1c
ZM+rxRa/ysWDxb4IyNmC5YTp81dbf/lGY2qLK7FSlQAUs2Rw8LZr4Qi2Pp8vTKsV2ym5BtcEdofx
OkmURhThplL4+Uu7y0nIxVJLAlZqSIb0RxELHV7qZ4L7OMUvgPqiFKFqMpKz2/Tp7ewep8joEx1w
iJzomAaiurs6IqwQOZgfKiOxu+1HFlwWgXCIKWlWGpOciRMFHlqwR/Hch1Q6sLRLtOsTL5wj5rzX
uoti1Q4RMLl+y9/FtJSxndQehjGqTI1yDBQzRtj7Y+HRkLNKkirjOw+66nYiLNbRLBielv4iPI/L
ta8ft3xJ2AVRERytIRb11DP1F45y/G5VlLMMtCmjLZH50LsivR3WZySFhHvIRmtkWN2Uw7L8Y/76
6ZI96hk/h8+Hd+ORe83HneMN7NFrO4VnDxuRV7cumkVAuBtqfOQJT3FiMzXnd6FMpL3j0GQ48ZPb
SqKi1lPiJrM4aPEHM6zVyFxXs4yhOb3YE/QeoZx2VyGj5Q7kYEHmxfAaBeQ1AodIJ3j0U2X3elBY
fMfmuKxYmxVG1dEx4Xy/zc4/NUSPuh+35w9mjfImWEAPeSTalB+XB92i3ALuuyzCVnHUb5bfSxyK
7WjHZVpVyituOrYd6boTgoudyOo+atwzoBDH+PqnJSOv4b0GxrLGoWuj4V193/IHrPeYO1vURZ4E
Sf3kE33taaIftBtFJyI0IRBXD1SvHV1nnupqIOspV3HdSaYtWoTRSHCwWoySFO3imXsZlleplDlV
+r60lb/PZsV8iA4avrqMVFQaNIK2yd2PA4JXkENw21HuyZjiJKvJlcJfUTyVE1ZWOUjMF/lW01IV
uZ8kBlEbf3Vno34yv90w+Imf8Hv8ooi0NEoNxAd/E53H2R1zWWmUZwF1da4d+kzfCtnPuWHtUoDE
z9BZZ4CmeYkEC/mhAOh63ISGdtUNdl3sZz8SMH1F1E134xirYIVT5Z1p+BqGkiXqCxdytZP8hGdz
AKoYMdgclxA17LT4AZLwG3BpE8unhWdSuOVSbcH2f0rThfRslFS/pTqEjnpWULoOgfhun5ipWCtb
MP4u4fznacBZopEde+8M2jiuW4nm/+1v34ZAVBMM1bR0grfNBvaUX/irb64pGx0g0bbrMOljCQxt
qU60aXj61hDdm3IW6qs3iM7mkqH03CESgf53S6v0eR4zet1T6nrTRPLVp8TXit3OeeAd6xM3ZRn+
W+z+dWypnYZFkwS+WJHO6TwNLyEmR5pQAOPrmA4A7gesC3diUZ7ZFQcrJPyL8algqiv71bt21Ej9
Bktr1jDcB61XufbupA6y9R2z/2Krwe3+RJjLdDgSqFywmsEqvof131LnOUsdkfV8Fc0nM61P4iM+
jfQsOpY1Ilqoy9a2pShMTuIH38OhEi1f81fZs85tNisdzCjGlejv4Nd9sngN5fyfuYciS4Ius2FM
MQGVUqvMkKk2mV/t6282cGC+inb6ikRIQ23XxDzcfQl0G7S365rqJUr4qLDjs5I934tQXGs5AItb
vcuFezGvsmfcWCY0PWtt9T8K7NHa0hm3aOYiM954u4iYXzjEgevzagz1t/qP3bKumdTLQE7AuhqH
J/JpM1oFXvdI8+mXUvk1uGSvLtwMsfAfMi/1XTFcFOH5RjA7QxrbPCDxyCt3+2sX1qswDI/At2Yu
ObrhCOayL5LdKgi1B/NsaCWRSBhGr60SHVoYXr/e8v1BWs1MGC0Csq2qxezqq5mKbDJFwkHQQq8U
orLraWBqIKLL1jsDO2Hbqa5A4GN6+TKLO6fjGZsk0VM0oekYKmZHk/i87Bhr8zl2siUS121vS668
rf8LD82PZQZOJniFTEh0KFct038OmBEMLDNjDZRZaUNBCyzZrLs19IsKMSzHouxnhbvYGqkfn89v
DGVTd6rti2gyeSZMQbvEgnAJKFGpBcdUMKyqHajsUjG2ircxXh5bJs82rlcQmRa6N6tWlQvnS8jj
nNz/csv2RvCc9fBK2pfwq5kQr10EKjWhyM+ly9DPh70gifpV3Hs1X7BSyojO00W+S6S1kIYMG5dx
dzRH4Fsmz4sAUSCPH4PKyLcn+uQTPDEE06DZFaYWsPiXJwXfPDgtLi8whgyi907NUKmLl0Qc3SM9
qqvCz7g+jc/iss+cQl0QCzBcyVihj5Iv4vHOdE5gfa/+bTzK5+YTtiUqf3GzWRQgVfiWVG0FLwDe
U3yiTXY48SOOjRZqIGnFtvQVlmmo0pnbNLdmVCkVG4TjFm2nMpuJ4XHf9XQDLLn3+qlcPkPVdw/f
MDWXe5AX0caN7OPDKb6RXswne5OKO2v5dqdfspZDF8x4c39QpFd17BV0QF/SqxvPGr+gE/4iBr80
Rf1ktgaTUOW2DLIJ2XybkaJp061dMqS2574dz1A2dj7pHPx4JysZ9s5G0Knz468BfoSXPHzZAn9K
TC1x8iMQ2LZqBzJMW59hSmryNjWHJIu/1t9ioD1QS7iLjYHkrOEO6UA8ie4DhWwDCB5xerPpIZpU
7FToCZC+dz8Mg44oGEojYC4SDzWdHvcwkv33pNecbYPj13d/Wgh1e/H7nYyJU8K1pupGTQhHf5wF
H/8rqXe7GSCpqbjobs2zH9s1DMMZ3WwhOCVrJiWfNCfa+WgT0G+VNp8hNYz4KZ0I2TJABdMMJq/g
aJgnwNvl5dHUEth0D3IOocyh4ymL27SE+v+ckxqjSdbLZS+ZsaPGTZ0A3Uu7TMhsJOWeW0/tBKtz
Yk/4hhrG8A4EDQcen6wVJNU1IN8issiYgo9dAwT+jisPHpzIQA4yG/kpDiAi/IIVdV0bpqr/2b3D
+2jgqPGNhKoy6vW2U64q4KDR08QDGU4DhZfU3v8c6l2TIh3j9yg1ot6mJBRl+3GVR9c3Zrl5rttg
7ASyVoFDg/8+OiuHC8zTENfQrt6ol5T6jDFNcQb0e7MThEZ+aQiCrXJSQXK4mQeWSMU6hQYkAvMo
txNI3vFyNFYbkg2oGbeDPuMGU7CogUJ6JRHkmkMpTtoR+M4/UkbymExAY2t2l6fVhVf1aL0NA/hP
fF5jqahzNYPdwcGaPMipOoqm87pgXMz27MnNYkYsorPXQbr0+0wRtDc90pmV7AVXJzc/ZMcPGo+E
Z144oAZn8RsHiNM9NUzuEPuWwHeuE22wJWWsleSkII9V8ISPUkvo/6ujDa/CeYooDWE4qt1amZbB
fZVg0zYl6rgPxAcov2JKf7fq5TBEwSLtBlRZrd7G/0V2XjthY/4A+4zXEvESI+q85W5DN5FcXJod
HDliDcCUUpaOk1wzpfh83LMQ1xefPbO1d3cjyDVi7y/jo4jKH8CKMWcL+Dymr4xgAnYfveiaTcCS
c7iyp7H85RtkpcTacQaSxKm7x2XrcbseDcBfilcM1lo2ogkR9B7mei/9AUj7JGiORhPn66fYLCUN
xPo+DtmEP5wbI68iYG7stksdgow+eT2AfiINVStGj5zP9g78Y6Cia2owN+yyDXOzE/Gdogdodw7F
vci7ckkMjQYcbEHCzT4vpJND1O3iGTuASwUpljPbkuZq9rkaHsr8AcBY82dpHonksAhpU+D/aVsJ
PfWWmHeaK3DevjPpXUxdMTmcOdBdeWX6LlpB8NHarI61ren7QP/h57TIXLKzrUCQZBfLRW5PUNos
PSq258x6iJfjRBAn3U/8t8kWKs/KgGceiReX6loXse51h4TX43ogU7ROaIGqe89RxrUe5VWCLYwb
7K79byI0y8shFOmL1u521t5mB1fuWJ89u13jS31chxFK+8TuCyW9PKXXf1WBCre4aLoCfN6ogHDf
7uIOuCR5C113rvg923uEcwwV7ZiZ8YKrsVTEGUcwTdFydbAApCDV0meXJXyXpF5PdQYltUeP9hyj
kxRg5oIglvx8WJsuONaT/vISeAMUQ4T+NWMcX6poLgQ4HzBfLX0g+NWOw1oJzxeUqZwK0EVC8eR6
OpLl5bt5Pi7I/cTLfNc1WUJ5YMhXCHarkIR7co8U9buPzhVT9NjeFUhVMjby5qExUI/04ktyNaDC
4yBRzo3CsY3IO9kv+RTJ0O+jMG/5KltvuVRi+WOX6pnElGKLn2vu+D/W85yHOxKq7lPllwT7SEy/
/Ijkmni5P4K8ngVsTmezsqNzyZUu4eh3a0yeGoB5Y0K+/e1XbN/WD04VG2t5wT3yR6t9L6DA0MTS
vqeauXtCdjZxJ3d1Kz600ER2ehY5kY9V5PgBhPG04UUtqduhPqL18y6KlBY4cUetda9ez19wNxTu
1cLIfuhm8s6F4RQJMo2fcKhKqlveCGFoP9XbWg/UmTH+o9Ki5lWpbsZip7D8KliM1Tx8HDGKemjF
QHU4x4+ZAQjiUJaNmaX7KRqJpO2Kti7oubAbaufS5k9vnB0pH3cjBbBB68WIVGqWuwsWU43w4S5v
mMTrFkoLloLaTT+47z1F4Czxltu3Pn7aROhOF85nOARC5JXic7wA1b+gLPjJ87eI6vN02YxXO39p
u3r1q6afSHEXcGWTf8d4RbxEpbkbcfUvfkIDTpmoz+LXZvs4vFBD3ghc8gQB9ke3kEwFLVGhpnS8
QwTqjlkAjMaZu/2bvnGEz82ajO3yvMs8AQXesW3Aolpz9CuWvddK90HRsgGOgRsoEg8fm+lI9ES3
IHgVDTBtRxSb4OjgzsSRnxXws2XFlmSx7BZwpwy2oLL7uCM5A6s8rt777N+5WbiU+DI7j7SzqsAI
ig4kOXv4dqx/WNkDRPF/35ba01dhm6eodyRx+JTeVHRhcRWg+OdwQ7GJ722u4POLx6m+E8G23OK9
g8baJQ2PhdcuExsnL5a6EeHyVllSFw11RCxd6tmTQ/g+6bA6zrafObjDvAtnqMvTizfgQjY01C+L
p8XyKmg5BzLK4srZTHAN81EMtRMn2IGF7g9pkf9xRInU+qCOABZbty6Vdb4lD6M+ACfecimjTLQb
mT7S8/r3sVF1ooI0YfFC85bGfyHeNUlYqqYJ+QUyYuNBby5GrQZn6wBOuU4gw0aMNMFEm9awgSQr
9s6TPcaK9p9qmNFrCvPS+ep7/eNNT6MYpsKd3IUnYvtZMMdNhBAYIMcGAFzsm57wqXTSwy/PYGsV
zrWM411YJlRVwpmi9/RTbWmUopWeAGz+h9m1suVO48PvQxNe9rPMJ9NXD4Y03Ee7cAnPThub+i5o
GGtK8iaIxFRxvVJz+5oFDVtnu5631yOaNagpxMexe5xdZnCppnc9trAYT7EUng9Jd/ILXJjnoemz
zhJPgbwGDyQtDGW4aHCE7vMHAzuzrNBtJWKagBlOn/kcnio54tcG3DcIqa6vjMbCJpTOdsxu4/HX
Y3fFJ4lxiQ+urLnHvB+Y0G3la7EcePqS8WMCaFZ4Cu3MgV0fABuuuYb5oKBxGLaruJsUt7JJ9lwM
X3il1NN4TMa/UuJLlUVV0APr57VXzL07tHNhgodFJtLzvlM6jms0P2qM984taQ0zwyyG6plLiGZ8
EZdt4XD+Zdt1YLIM9SiZrlAbaxLzViL7xjLHppkjFqSmJ004ak+w5+Iyij7eVoSLN79UvMc7yIlu
P6c3WoBFcZXesytrB0HS8X5sOTj7mzlrXauHzwp0lgFixf6SHmnI3aIycSuhPNDXY5XG9tZhyGhC
GGzFnhtfMoJrBxpZt7GjpWk8v3f4UHV4taasRQpOCiNCN+qjQbEyfW6gok/Ekw+1+YsqfT5krw8K
cQNctp4Sb2NNRZY/fZLk9MuQPZgnadP9AWqnk14hvCNrj3uEGBPoJn0/q/9PSd4s/3HdSWGkuuf8
2A71rP0NUItnze7fPDCI0YUW8ddQEmo9s7KA/RGJ5d6aeNofnnzOB29zOENo1RnodBLKjLsU9lu1
FKu11nRKIX0neBsfwvdjaGBBIxItwBprqC2r34cvupQt7ZUrbSWDTEx3JbnbbtFUtngPk2pOCqhw
0/ItC5Z6tEtgc3o+U6aL5hAOpencqUgDI2M5q9HaHYtBEtcySf6LYl6MoF91czG37QRh9e3p1ad3
OgqRkraJvj9dsPwICTW2IF+NGjm9awbQImqKFtd5W7OqXucZVnNjm48Kz18dMuE+3Dg3S9Nb6Mti
uH3AYfaBkSlABwnOu/qQZcJ4uZuq9LhgtybbsEKIg2obv+DCT8A3FR2TM8YeeThURAanRUUcQPwB
Df7wWykpwa1hj7r5jTLjL/nnzPMsil+JObaxMpt0TqCJsQqVPbmi//r23M61f8TwexwzotHnks5P
C8XlGLFLpc6whVPFiGaaTjtSmVyluHG964bukaGp/r6hWlEDtZZFhMTXCMmweElb0Vf2Wu8QY9A6
6aO64J1xDgwmlDsp3kAyfzAcOXsZtsXOwfK1m6GC2rS7NwiBaHej8F7YAPRNLZCqxI7AvS0dsIqB
iJvn4Yn8O8bL5tCDrzy2ltYjUnyU+iWBJXxtsmAcRroPjG7KcE56TliqHUt0G92Tc9eBSvlBBjvx
INK9xwpb1cOBRFOYNer/L3S33PZFNXPJOvpbTf2syFEHvKSWFCGzus8wKTPm//LgJzXauGj0nrp/
miK6OkoPcvjnkpQpG9h70T0xss3wTDfXL/9lfmgjwSSvabVKvqh7s6R6egNe8uSsRe0rnJDXG7nv
SgiJK3w2plr2U5FoV954rhWIcbPZYeC1UZ1Lu4SnQRXZn//GBF0dRBrTwfoOGeORcXZV6IyEFU9z
7+Y+XiqpDp/6Jmx1LR11e2/X++FLu0spu1LH6BZFoa9xumcBWyzDsGd9QXK9X+k0tNmkjyo9Sogd
SVhGHDyoC9gOFxHQYT11WnNL+bUzLoKWNIxXtoy16PsXgqYTGYnnRqU0Omaej125bGDpEXc9DSx0
Z7IRX6PX2p48m4hkJ24mMhyZCoeGdtP4Y5t8of7KjnpVKOPe0D0ss8q3xwFVzeTSwoJaI+GuovaZ
VReZv2dJ6/aeHPuSEJ4BeWFFLXgbOG6kTsEJtFzG28qn+RZZCBERT6FGiHaNaYFeG4RpQOv4xmuV
T+VzZTaXbcKCD7AC5a/kNcXHnKbPvwUeuqd+95yoCj63VxygXmXlTch57KYE7cT6sLS8DT+yiQZ2
LTzwY1ouJOINPGj49Oej66Suhx0FpRt86JUQU1OwmgkW0nA6qvPzLYmtQhgaDgVHic1oA1n1ViAf
JjEmfjmobHKRVRFSiIAwUbtB2PYRVy1UgBPr6XFivifyZxYHXhoAuG4cnDi2HT7MN0EfagUOO4Vl
qHcI7OhPgE+8llVS6npIRpd8i2GKyYHClYQM63RfFH0eFe9Ia2VFulHBg5DdfVI4qZmGALUpH0H/
dMwc6/bpj3x9OArnbRmqh6EjO789bzNzM3Flzj3ZYGhq8x2uOZRzi9ZR93m9wWVGOk5gU8/ibuo0
9cA1qHkjfRT+AY8QQN7jkLlgNthBH6xVTnLJaKI6eF0cuq+qE74trWMDD2r3VwZNRgTjbHTxZTxP
3uoosE5ejQWMvWkD4yjtfHrRVWz6Aw3uTM4CPa/0vMKe10aS0EgMJ6cnaPRK2FzLBL8Vh4kuTGF4
Dpz9k9JpRKv0q5exrT+fFrUbY8uF0uOff5CPIG+hgOguwq9mTtEj4pyrpYEwIvAiVM5vrPwzj1xA
oO6MiIRMdW+3I/NntuC/xgHNEkI4YbIkmQpVXV8SWo2XSPPDOxp4eZcbSwR/ajWoSL7hVM9DmkzU
53epePVIuPjjKBMaCscvPYy0gRQae8Z8zF4jPX5aa8vGt03iwWhfuNf0CsTfezq/mqqRuDLAMyps
Eufc0HA7Uccw+RokS9gGxR5Elaki0rjfd3HHPx4BwM/K4ZMSwM17w3DqayOID7RogJqLeUimxGtF
3dFs2HuVX/T0ajej9CZJJWIgszEp5Sqw5p00jeVBtnI/cJsO3Fpz1rok4pF54X+Ha4vkja7crRyM
bXa+kaUJVyZ6lokynUM0vscCXUNwgwLt0FDafANjcK3ncVmp59o8t7tBv2s432z32fjtFXCqbQBs
ziyFoGj79p+kuIcaCETxKNMfCQCDJbYXzF+/s99kfnQa/36myNgTb8cLgAjNAxQ5GE3ubD0zlTV6
VR0dAqu8tzNv583OfkWLxeoFZrNVyPy6y4OupeJ+aP4SmPoaK5DNy6lEt30bOhX+gIMq3ZPpnaGA
VGDSxUJ8zbawyFFNf5pxHSAj450jrWr1FRtJ+aHM1hu8Vq9eVBQ/XvWva+Z1YWKQ8yLeKwXNI51k
3QJfonEMMF8ShC7pFC/0d2XX5xGB5fs9cH8u4OsrvHaoacQ5tCQJdvMh4XDSK75mNkahjzbM7gGA
pZNcoTP7rdd+2o2EPhNF97F8b47Iqu5lXR+hvP4dIqftzYbsrWzezZoZM333ikO7Fex6tvTdsMkg
s3LBNrAoeekiqVdeisBPdBvmyrrSRi66w7fk64reDvVDYb5wPxynq+XNtw1TiXFONI8cDjW0fTVO
n27c/BGLYAZjx1CINPHBzTkMd73mWk7b9Ik6WHUXENk2zstsXfd4Ds6LAYBQZRu4z8NIPvEydxNy
8E0l/jtWVzoq/vYl7IdfGMvj2ZK5CCwdEtqJ93ogdkgcjwDcHrKm7cekb8lVTaN2J2U2gSt5DKKF
A1ufd6Ld4wxfI/1CJkdgKbrIPB0MIysaNflKtQuJNKUtHlZAQxl2DRRee7+zVRBrJkTSDGNfs1js
6pxUlKxYbJNLIeRSiNNaHfwO45+bB5I5x/c7sHZNH9kvJuVHT7+RftuaGMUcd2uX0Z6zTcQHXBu9
GtiWzeHiaKiuuvDbdjrbwXzTMamXSV62pMwwAJgujFFw58n/5GzdxlydC9oE/faQ134nBIEqm0BG
BWz7BaqfWf2F1iuxSNmeC8untkia7Cc/kO6il2UqBqQjmG7Jdc3JOyMRK4Td4WgxViw73Lp33fSl
TMCefDkhueOri91ymlTvz91Zett9DzAcbAgpuKB4UEq3KM9CY+JrLrc48QkDiWpvd3JMDocbQ8GP
zRGyk01n6FiGUVz10yGkNN6kyzxKVB2RH/VKfwgEZSJDfXxh600aQUl5xjmHVAWULQ+w88gAfv3I
eQoiaisHuzHcvG2cOhxSOH9GGEBPyq/RSUw6J46xKu2D9LzlwYQzFpfCgXklqX8pB6ZakTYZjQUh
zA0eBu4jJCBZWhmXqa4bsjExVIwNWTRUlA6nCVkR6rO0meHy+EuUN338cj5CtkUs/FdPnXkPX0YF
iAQXA0XxTf2slvAS8IeMpS0W8J24M2wXa8oP1OHB6b2DIw3cQjuA55wqgn5NkOm0yIC+hsDMQxWE
oTIpH0smLJIXfyGrbJES4QQoIbQYgnqNowlJMdzphumSrSyvBjJYxP7idG8equKMafCCasFaA0dv
36vHZ9nIIdmhHKYeJAMo6k7p8OdS7s2wYVc68ipF06VN6U/tOSa+au5TCSVeJHm4ImZ1pMkwZ1oF
pL7X41dCse/7qW/rnGhamDjZA1vQ6UOx7CU9ns5Gs8SMk+kFx7n0KvIN7pHcq046YsjGM5LCA6B4
Tj40NnLxu7YZ9+qhB6wIt6q9UN6iSUrp7A+W9MLvMUTxJKnAxeQHr6j3IDQ0veMAzTUSuODQuknq
xxC1JGdIxhtgix1N0IaXeNVBMU50Qef/benUIylBZz8d1Afy2M82WOMIuWV2vHMHpVlKPCmo9Xan
laz4BsrYLtA9zU8EjrIfTdvtmDtJg2fI2pH64OsKg9hn6ziILCx9pbz82ibOA8NDvzt+fi6340hm
5zy87K6H85I8Yakfz8peXj10vniPwOiMTWgFpb5W8JbE5b/Z3fz1OIIX3SgjQliChKi+zjQrIhZ3
DYFqiuR7JP4De/Qxw5aUpy0LxMtcJFasYL3SOJU2vCwihcl3XRMVizE+wjoBbL8/CjtHOlwNlVfW
RXvtrGcLWG5yWzUjckx7ObMzRf1C/t5ghAJ/qmtqwDYAFTs5JQu5VmclWUuxjHid5yMnyPq94tZ6
qyxEP3sFyfM5D/sAZac57KngWaOh4+EQitfUjfok5WVrpa0OxIw0K6SbAe5fjZEHw5pskBSF14Lf
ohWDmzj16STR9uQ712dv1YertcfraNhDMVLy7HMrpd80wQAtVLBHTfn8qsciuHyzjE/kY/8PXgmK
9JXH5eK/juZw6rQ/1tmRvldy+4y+2+kIHeMGjfZ1oJphHxi+XK74YYgZX3X24fI4g39SuB7BVP8S
8Rk5gwZBZHhbT9tnRUmUr1rOQ0jPdYiNbXNRtYLmo9Tbtw3AyzK6n2Vm8ZfVgms1qJWCEztnH7FT
bYZ2k2wswjgOrOjlSA7qt8l+zUAI+gsG/+Qg/ud086PNhkCMhCm+UWDfLYbGrcbb9YAbegpNbHBf
MyI0dmmbuh7gmjN4w/7k/MAbY8CjJFxXPgJYabtBRd1ogDIbszATnwZ2nF5daVXWBYPG5I61pfqk
cc7yuDW8YkBg6Oc8SXUMEPHO3BsisbqhJj/4dyh5LQoO6yzg/7bHFBP6XEHAJxXdByXA89V38OSn
T7qlY7Kca5Qh7JKlq7C5erKruRKxrBnluix5Hrt5TfBMT7xlQl1XNZW1ev7afhbnTjHqu67q9p0r
H8PbCA8zXrz1VZeIZ2dj8Ne4RoZG4xDmrYUWUv899Z9W8dcy2el3bKsHZ7yQctNELNh8z9RYWlr7
NLoqQU5CxibTu91Kew3b0BK22DvsGgalSIHB1w6BvCOKlHKKGTSq7tYi0/Kl1k5OkccVhG21HtqH
ym56JLVDyztbcgTMYck/dXvJ5nYVvquNQyzlwCitJMEkpk3TijxQzrAmchtENTux8Xn6Z88TDx3P
9M6e0ST71uCmGLWHcoK5Sh6Zh2w+kyKD9VHc4kmENDIGNweqsOPPsJ6z4lHK4ql9LJxr10ruv+uY
5H7LXnxmK0c2Kvew+BzLdXGIPMv2Psd+/pTbfJjd5cgMn+TUHQM4rxEKd3jtOY3JQeV7g0GIbQtg
wUAOE38SITNxlLs6g0o69rON2qJW1UMef6G+jqBokOWdSN2XkiJr/BC6eOqfmplXJXWebTjQd3m+
/ZENF3nGObdzwK/pUF4AJVVOvbbGYd9OecsEW3vt0R0W6eWQeBCtKGxS8scdbukMnvpVF4lcDA0y
MAxAbrp6x3f0asM830/xeQ4CUDtH2Xj7i3i+PJKgsPimR0fKBgeP/OD1YWNzVBV4miRvljqLDbwX
iCyU+psqkxptAmbXmkfWmB+2e96jSmVvCQyNDPH3Sz7esgTrSv2bF6LDKmVadHMNEqGb5XwIt7F+
biGRS3ZADmR6KdLMgp49uVy/KUAgK+G7aZlsL4cKof5EeDLLtH5DiFTiqZ5bIITu9tj48P4jylg/
2fVv+J/Xllu3ez3koZwVsL/9WZBGT2KFb4zZi64CNV7IucJE9NPDTvK9xmldw821tsmBL1G2g8EF
7frb/LS7RrAuFvqPf8HVZ7f8wcXuc0LEUHXnbN3DYfRJd5qKzRgvhu7paz1WBmov1eMBYTH6adV0
g/eV2m/1gMfyW4+J5vayVQ0M4Dt5td+LxzsRLPA1+zqrxp0wxxzjwe8rebWhvDUGxkTu3HFzRgLF
wIFpkMtGspEDE05Qr2adaCqKSeFTGgFyVYm/d8hYTWVDfhh045J49g6mSqem2C0IoUi2Z2Rn6FbW
ZIS0LGtAoqBEpxOgfqybn3fkSEFjTvvgHMmvL0lEMuFmN19Qg4mTPQG+zHLRE9AD8hPbsgfx+2Qu
tqp/Gebg4OECEQnuPNNm5slsPtKimp9mt6YDbl9K6OfUgaKyWZ+zedBa9QpdRjkqCu7x5RPOwhdr
vcacUgud7UgUVYd8q3tsi+wm4zEZjhgOaPqDIdbXxyt39THNFexb11izNC6DAnU+OCsYtER829kv
R+t5JlOwLX720dzvfcbHKkyJRZALC1AVU2NQbrt3RvYsN0VWFZAUuno01C2Em3J2W+XTcZM5WOAW
R4b1gmSkYb/ZLnhWcOkg3+Pxsg5YQseXqrhg+HlnOZfR9g+p4eNzf8WAH5707aLmjkNA/t8DFb7+
HTgQVA5r+yspc4F3VU0mSsTWkd2aWD5knWFyTlP3XkUlK+L65looBxOEuO5csndmRSh7dONGfAce
dA3ke1mRXkM2A9ydrZMyz4uqMWpbnNrau86zRLgWj02ogUomkwbbSwRAJKvWxuOkkI3917YPSr2G
9Arxnla8Pq0MqJ+bVvOSZGPgMty0cyKrAklOOKtB9WxmPSygpx5Lnrk+j0yHNUNjhW1Y9B2Dao19
GLADd7nn2mhSUiVQj8kHurW3sz+H0KD+cvrV8oup5E8VjrOd/G7x+bHl5mQBvFNXeTI8xV4l6pNq
T2xW2jaiSQCu0/VzN+Stoda3Dtf4rnz/wCj/nr3MSQsqtg5bFWvS7UoNEehA7+YKqnPQRRApKhOP
Z3S5sJKUa5AxdmbyZAI8v228VwRF9pWP0nKFSTViSPB2K3g3UUSGCxdxMlM7pgnbpf9UoU574tgK
n5zzXgjciDahgkVxxUesk5tPnGujJ+wMNfd/su6c41TX0aTfz0S2Gn5YVwpvYxl8p34L+/bXHBqL
m8ZsJjtKfT/Z+dc7A9UAfBvFAVIGdLIgQJSHmF+nLOZQuKmbgWaP5wSMj5K2mjbtU9z82G8zy1Ym
Dv1pR/V46X9bIMPNye0+vdvXtuWPRMDRDAG78vuSnx3UB/8dS0otPzPCLyTKpaM0SNzmeNZjyzeQ
boap1UfS6ga5IJnRXJJ13KKMGD6G1LE03kw6itmbCV5MDKn2HBn7pmRHYxQFn5MHuIGAo0zsSERO
UmtjsJmp8FYBLWuUVtan9MAgdYb8q9IoxU7vEqkdgELwqwQk9tQsJWGf5DoddCgXlQc/g2oQ3fA5
DOkrmvHmcFiaLY8Lvu7WCjudD49cqB6SFpKXwm2mOaqiAHcv5NcxWGmdMj1zSqs2+dm2L6dL8ylR
oZz69WZKtiW9PDuj9hjSW5krWXY6zNxMvFB6YV3qhdH1YYZHJcoerWnN0HaVG7KlJR89iC096lgd
AjkxOL8jtzzRpGbeHmFMM8MaBU+ESYKlWBo7Lks3G+7v/rPsulLvorXQFz/ZtEiOCf8gG6zmYa/R
koyZFEuIyxeswwm4NAOQdjv4mwouq3H8ek5t7h0TmkHLqM7rluk5zc67W+0taytBZxrR0l462Yvd
e9xx/9BQuIxvsiTFh4xKQAInPpy+0g+ls8MI1kQ1zq1Nyy85LeS0qga2K42A2SjysbloBiSPj2e9
vYhjUMR5yJypt//L/EWW3AS3TIcMoKWjKQQcWzrRQ+z8XBv8fbeV9ggFtZQ17QxzBhczxYXMs2bv
iPiFJMAIHaFrVXi6BAcd/+37LsGYk6hTF4H3FOYll0FJW50w9q3RM+8ytQ3g+L8G6JWCrh4IRT+3
uIekivJFtlucejpeSVL6gtiQ+cOX1bTOH1yaOt3In9Zjtt1PFiMccyJFm0RWMAjW0qG7yRuQSY1+
jjiC8XTXNoNKE7afbbEtp2OVSBNShyKtiMD3wwMA0Nr5KZKmGDRgS2/iMVgb0+QhNWip6Xoc4b23
5FB2eZsq+OOJrwl2wOkNdzJl6QlXvToIwlRPH82w5UtmpQdRgkizoFyDJZaQmognOSMwPqWLzqpH
ZDHrnsC7cQB9YLl7JzaaT0v2ulIXiwXpR4BvtaXHpqY7gpLDO+Ba3JP7b//pzyvPBmXBwX+64eG2
BZHfNZfHpXmimhDnNbVVLg40r8d0uO19+ZXoGD/HcBB8RPg3E4Umrh7f6nA6ClY/5A6d73t8o/T+
sFTdM+V0oZuEoFyQzd4hfGosTt3KC9O8XsWpguFUMacHWqQaMrii+6E+1bW01RSoV+ZA8OZ8EKMg
eTSmoLng4x8n46YwL7Wy0RAHy/VEQOPapBc4B/IZdw4WQbx6aZwunOXlYwE0geguB7DUCrx0EM5x
e+IpbZpMnOsLSysUhXh7BxASTN0qmq4VJbXNDKDpUc7W/uhuWha+MRrgWYXM682otLI5Rc/Iigp3
9UVBEBDySIounOiMizMr4st6s9EHubf6MchlR2O3QdXHEyKMhLhn8qOtB53LMFE6EgBQjFT+HUHJ
IFeFK+A7yvUidh3RLCojm/EDLIWjgrrD+BqgRU1EEWw1QJCM/ADQOQQ1mr+6v1tDLD7z1g0cIFM5
wEz04pJi2GHB/+eBEFoa8HH/KtBJ8Hflm+TAtjZD6k6C6RBStu+ReDRhD1RbPseKV2mE2gtsvK4P
3lLmKbqiOmnTsP4j6ecS1iD7qe0YrhAn/Wpw8nKI0e6pkgX7v5+qnOXhe6JMb2dkEiTd/XHk71IC
Zk8C6cQSKeEIHu86szGKPAa07ER53gpl7CE+8tRl9wO2ZnruKYgGLyVimEzM96WrzgWuvFBAGoaN
dUeUrFH4+7MfKt3/VhX24Gcx8u4PZP4C1HiaSjBne4efv+lrWZdHhozXO2RKrB7RwXpE9DFiXHFy
LY58esoXE9rKTTz2GK1YKWvyBXiYeYdBA+QEMlqx8McA21g+G2MvPVCsrTMFvJ5HCGIyDWEOk7Ww
FbLbajoukizrhrSwsmgF4ffZIzsqF8CLMaSztP31ug/vA+0l4rGcME2A0OsMehhl7RFQpjROn3Ml
l5D4UZ3t2zyAHRmEymusZ6aXfonnacbQ+assoU/Y8EeEIa3ijyhsz9zh1HxU2kzByH6IQLf+0CLn
Qp5KUYk2Re7tL9EC00fVtNyP0Px297dbMI1yTCMpucWCm2NaPUC0ts1vcZQ7aU7oy98UpyPChGPo
TKGmgv8pogOyTrlWHBTA03VlQ3kOySuo0BWV854fR32xKDhbdElaNhL1A8i+rpGeJWKm4/slQKkw
fjbBU7sxhrkXEcYH+sc74Y0PHCJMhspZrR2FSeNlkn5oh8ShREbgquYFm6dhSIQuPYoh/0eGbxZb
giePlpXOGjhdUwgR82/wyO/3xwP7a19qFEr8kDC08DCV15NMd9StLAmIR5rxcWPNIgipPi/N5Tj+
KVJGmoUSZraOQC57PB8eBXZYGFgODWbrD3tkLGgAtfG8DS1PhbN/JpE3gJD0ee55ITduOmQ5V0O7
JmIKsx3sxZFdJI+6bLe2YfQ/hxJ+7ujJwEYJn2tb8JPdKJ8aQ1GvOQSfER851emPTprNwE/t7vcH
hsHCSbDsCS2eFitUtuWwsHmPIxs/L4w2wEb86UnpeJbXO/kuS39nHJqWKVazQuwiCdO8OfFnvxr+
EeRJTrr/fOXjLJP++wk2nas4+Yp7s3ETfzAub54NYcNCkIAMTb/Tvci5ckclSF8ch8vlU+XjEooz
HmNTkFS9cF/z37vV6RilWD2VB76xaDnp6yNahk3EjoBCz+/JKFus7yXsV817axN9aOvlS23zrNdS
LJCvOoa9+JevMcmT05Q7KNM6HMh5e1DdWbEEB8gU+TTV1ytyMAlqX+rtQtOpygfcNPuf7OaJVIjf
5i+pB2EoI5gApr0W8PdQtsmtOQOVs8nPVW9wZONDmNLe0AL+SwRSPLFNp8C/9oDvqkx4BGzAGRDk
7uTipwSdCNSDPb2+qOocG3YrKwEnsNtLRPkvBfuYZJLs4oQhkqpc9BtJ9Vgy949OYD9lk8HySxRA
JyuXx13xB2/fibpIwg4zTeisMl9wU5vgOU3M1FzoiMcq7RMoz2CnpFDsJS/oe+basgIvgYkjMe0B
8qfTBM8XvCXRsMSh35rNyggK+7y8MQXIafaJWqnfJxbOckmJanJLTLdUeVa4xMr9W0xswJ/BW1+Z
I2VzLJscHLswm26rkFxCdwOUCN3ZXklMS2Ls8UWIiwbh7pkiEnvaPQnNc9WlaojimArvwQjfDTPb
M420KuEC6LMHE5ABtLELrLwZmCw/QCf2YJgN8xVKduXV9bBIydHqnt/Qy3tR3b/pK7/ycO3HBVwQ
p5RURGDwWbNmGQQNA31RliDwZ7Ez/acM/I1WV+HoMrHzAo3sEdIzZLBRZUMjLOv7wuWjp0+GttZD
k1jgyvSwRprkZJ45jiDFrPoLXFt3DMk0r+GA3wBV/hHpR1a+HPIQixLgpTMXLWVxYuVNmMjyg36z
CVkefeJUDvsFgRh1CxomL1l28YEPB91IE7tfOi4gpeaR3t+tzN8BQjkfokqV+KD08qusPbn9f7MI
2SU+VKscunx2EuV5/3R6N0kVYKQlvZP8Gn3iG2cjKZcIBwvFBbBy3odE5y3ux5jLgTR4IM+PHiOv
/j2g2JKImHDNDRzlLUdN+9xDgZay1gEzJvUpA4ioUoS3oJkZBy0XVO9IqXLZsZHx2yFv+FffoKl3
miD/wMUsDtE+7KukrjXKeBzyuXZQSBv5jkKAVkKALEet4dW65ozhsLZ8ya/FY7sxX+QOGy7AFqcG
tedIoZMr89fMqFK6GUipVd2J/bGAN1t4wOkgSE6UsjPF/uGzbKPs/eInGDnkk1lWNWupyRiulQ0s
SzU4kJb5gCxrnLXxj2AfUVqzEKleQ9Jcbpk0dxMUIS3OwxMHIHwkEcSqMCTl+M0If/LDYOcmV2u/
XnCY1cTjDU/mjiMleMv+5t7nvNiPmEBBBHgjP3nlBCugFSQCL878lPAr/oDp13qZ1H46qjx2o95t
G3Y9h4q6eTtITvHNxFhWjgGr/Nq3dCo8JK13bBOz+hgzopAw61XJB8lucO+Az9F7LraYnLMELMJt
plv8hr4Y8hcvh28a8WoOyok6YaMpMzGTcZTPQFj6E9GmBldzAJxXiM8hN/j/qbHR2DeJd9j6gKJI
f9oOR/ThaI/SGtR9jgz2koo5Fi0fT+kzSHIzj13Gxa7eAvbBBpzsk8AYWylC/YBgVagbrfZwFNSi
HmjbOs5aZ6W8cM1UhhMP9eRJiAhnwx+RBuPkh6+BOMWMoBXCw+umGWdHQtNFwuXqN4RpTFXGXHA8
+JhmFsM6JWYwqQndJJra03twVdQeBpgcQi9JI7MUGHv5fVrWOPd/W/W741ezkM0Z9BxdK5nhIkRI
lNOQ9iOFTKZPCZqSYonh3A1dvly1fXEgQZsUv4d+ourdkr/pt9LliP6bspqrgDUYUI8O2y52iaDa
yCL5dpnjg6+ccS2//tPFrotpWE6khLns3A9oAYRFcwFda5gxq4Qm2e5IrteVAYW6k9aQlcCZ2Lj1
K9Vf5LKN2Jt8+D7z2Fzd8+6gDm5v3Ac5b1aOITuSQJaGfXiMAbSP7EpZ6vNUqGGLUhqJqV9+fnqa
Zw/+WNlNfjCy0tfx4IwdzJ71zpf8gWZYPvd6b/jfy7O45Rp7byAwrPMPw+WA0JNSFun16lixCuN4
r6klWRk+6NuXcEEd6mejCuOuqEK/x7rThv/+aR6z7wMSGrM1TBquk+5XkhQosGl02pWkqoGmWMB0
TwLHkrQPefkVHIWPEBOnXkpGYBIiUCKr3DAWjozkg0keiBuFpzi3d//Du/O6DwJ6VrE2L8Oj8rgl
gux2qJIIXA7B4zcgfjUrhAeiHYKgyEZhymS98BK38NKAZr75SaYVdWTwCxLvY8MwsFFMukN8A/CN
dL9TUcflYCOnVJZ7IJH8MuBJ8dZZgT/so/87TuEcah6MslJM+DTEj9Fx8lD/Dc69Opynxqa+Rncl
BjyBS+OXcbaVC8nVDaFfEbFzzNlkMEGY9nTyvpQ8RD4gM5FcXjmsURs09uqOktIl/RRCBTaMVJPK
BrhIWydqVO7yaFrCpqn2WD7PhtESitWMk31nAYaIn48vRL0Mb6r55nH8e0zWy0yGzHI2Zt+cho6p
nkkoj1iUW+2qfeZbVbi1iBTkuHTmi5yydQzns00HdO4JwntiEvYHsHOyUI3Q9VTrq13ARVtX9APg
CWJK/J7Cnt5I9dotuhl9H9Pvn+JshbC8xMN1NMuOLVkbT1GZ91GstMlk6gnxiIsoEjrkBHzWpsMC
lSpC3OYdYAv4WxOKh/ZbuS5wtECuJQ001BeYIy5na8z+tdbAPwMbTqZdPy4TR5iNrr7FVD+9EQsG
BQUXWHl/pFiOTgP8Qex8AuvERgntreA71euPFqTgIHVQFHpqCZqWBQ7NMyv5CgjaEm4+mwvy+ysC
kz4ahBZnMljZmMZJbQwtCAq/QaipIIAvnIHP6g+K1tCwo5vsugVE0V6WNaOnKCNYKJzfiNyOcGA4
1W4ZPczX76RpXbQ5dOV0dS/q5gpcLeJGJEHy/hW2t0ohY1+CUhiTnrcPm/QEEflxjDFWtuTov6W4
ZqoyLLjVu2dysaEz5wwWihE8S8Ue+6o66aI+1qDwXA7R2EvboK0x964sgoeLwxYB8fD+PLR00OEo
gAAr9CwOHomMVgKoLt/m79oo6tiFZvOD6tkV+QeD3t0wZygV9x3bnczurH1Ccy6W4bicktdF6mWI
Y3Aw2knONcWyyrlembMc6u0bSMkPBLYLx7kOKZAg10dUlHlt/kxJLwSVurfccFfC4OaxIs1LpZFy
SwjSnI5izHAVKgPmuyUwi8zVK6OmSMm0Hsuh//hGo1N4l16yoH5bVPxz+T5IvX5piykyFE0Gw/gX
FNHunffN6Gtg+65byj85vmQ+O5riczMCX7N0kcbJsO/AMuyqJ6/JZTo+/taTgGDaNiwO1rXAPC3/
13J26GNr/dU5ZLYniQ4SFsm1O32AoD91A00p9M3T+vP3+BPvEtge8UUMAP3vEaKGnh14RslwV6fc
oF/eKhDmwbs9PPwG93LgPqhWjQ2/2127jYrjOd9EIUV+DJvCUa2MlOCQYWu+wTBSlEQW0FskDT85
23MnKQjndbW+lHVXLq4DcVeI3DE0Q/Xgz0Q2Bwpa1s0AUmO05jNTcgtuulRh3GqZfsCfw5ljMeRh
rKMXfJvmHuAF39GwP0JKGwimat9eUJ4iyQfD6GJHg2iWQwzyobaYeBWbkCWomNMPX+tV3l+hTqMK
H4ry00pIq9XAcG1KgXiyRNWR+r2R/KcSKrX17IjYPncra132iGWmLLIcI+3ptADEPw3tpAVcyrHe
AF5eqxnUOSnoRxu9zvNXuu3VigTLZxedNVknM9YJJpfVdWGoCrGd69cUNmZjPZet5IXNCF/JDKAd
aDgN+TVwfJQ4+PnDlGjcQICCAvwxYPmQQf1uaGJqP/7xkQAKj5uQWCSabuNO1xXgXC96ocnTejO2
A17vV+mlBZB/+he+dt7K/LckJkxT2lFU6d9+pb6VHzERyjEW0NwshFYTcx8aoT54AxOwFluVObja
HzWvD6v0dCFLmOnKjjKJfx+pFyQ8lDWFEsKDIttMH3JXozxQJtwp8VjqzTrYCTugu6aJcv9P7WG7
Q9OLiIVwAr/QdeyCGROaoXKIp+Ye336Hxizc59s2s/nT3qM5RFL5aXJQXE4KLwn7oieemVDgRAy4
EPc/Ii2C2s5gwfm1XXsz3Wmq+P/bQ1xq/DttBcIXkxMHMM3lvQx/E4XL2zBYVjH6g7yX4v/kwoIq
Vbm+oKoceOFW1ImINIrJM/Rs057NLB0fa1jk9XS10lz0Ne5Ua2TXXWBLeksFn+g7tVDHJzgCuQj0
WdZFeHNYfN+TqsZl/LaIqy1ClT3WcRFw9rR7E/EGCun+IL+CIC07LhxTgQ6SzmG5MRoAH803sjbl
MMVDTaHKGxyc69f+SLS5z72FGY9HUU1RkK0Gb5p3K14GrfI8vs+VFmLKtZJI9+qUEiFZGByi3Aj/
r2FE9d7Qk6uWzwMzhldqQdg8jS0l1qHyLLmt2ARVip13TWEz1T4SIiET+MbEK1fszCulvG6jiVA8
zBhjpZjBKnuGoKzBW0j/I3oh1iGz2CvJA6eflS4jd56cZVGgcj1HstxGlxgFrkPnHpYZ0zHZD6KM
t/uVtLjP8Ell7XWREEfzBVl+XK1YVEmZW39NGpmNo0G6f7/g6JP/Kh8BJmkT7bzvKwRmKpNasrmg
vCYnlcpbwYXuu2nlcVsjyT3KBzCECDwwA3kvkkRQ2Ms1E4x2jA1TN4onHXpFHrSfYseu5853Gtwi
k/AGMJ8/4xmuikHjS/T2Rl81FSxbesdh6ada6vCk+k5ydQgBnqT0fFaTmB/aOjbDdkS0EIqFmz9H
5XiAwZ0V+vUxREVn3y/ezBFSpxGEdoQ3IF4WbUXXO9siBFBZft8Qc/h86/U6Mb9keWzJlaulWBDj
XWo4cORfonRazwHkxI0XnACP2vOuXwIzIoXCIxZDAnIL90MjeU8PvuBKl8/ZKV+1eddQoWcm76/S
GgIFB5eOGFsVB7hKK88/SV7SRxVPDTCfXz6RJqL0+uN4jl+1TP5Xzg25FXvockU1VirJzblZb9Hc
dxdXGJpKS1m/4Csg6Lft8JSD4qKL2kGGtPTQWXIy9zVjBPvLUKsWCB0jIWhY2QQk1Kcchc9cWPOZ
PGMS/YrvcqTyF0h8DEggyYyv+LGALpRcqdspRhxmTCVfKM3wlQHP8jGxXmxJyD5ejcVutYDboIGo
6PO9Oiuxmrz0Gtv7iOUHF6djs2ygwkH3WL1O7fxto92mzBbcGAL4GVutR4gKxiLcYYl9E/1mFqXN
n5TyQGKS028ZvkSgFWKS1d7irqAh8GqhLP6NDWZAYW/USDoLTdsKh/psMGoFy7I79xOCAMJgmnOU
6XtS6aA5KyM/s+cKHc+2LWf2PgIUaOzuYcN5/Z+xGiHiyMm22dhtKMYcGo7yufCjM78Gwwzds27v
1StmoPkLLtCHVCtwod+Enzc+oSK8AoDTy+VAVBqpWx9+WFI2c2LC+Bs4JyIrl88kNksN8Nuy+gY2
gWgrjaiXqQbwKfuiO0HJ+rjJo7Jxz9gpr2f/aHIPpS3llIGpTMruGYzUQ4XoIE2UKLyIdgUNlznR
YBMPiBgdN3ZnyzRmqCCWTi+Vhqsf9OfQsqJt2qrkMp/6Aq2tKJImZug/eIzFh7Y6kcXD464ug2yo
UNRQXIr269mImLCHVrcuYA+Utyy4IsTifd8aaHm0rOkIfvvROzhQSyorfUrq2DYYvNSuFPm3oBtt
kSfjBPXC4oTGdqmpMstjTpmYrtBlpHnYI57x7KwftKsodpdPtnSwzUaUIKdh7olOUMC7lNH5MCJk
ivev5WWQReN3dNmUXCgMXAFY4ZgH0x5kFtm9god9iOoHRQJ4ybbWaJY3c0LcqsFKqCO+Nr9hH7V2
Z8UuPJ/0nL5b4OueXwp6oHrTBAXJn64EIAWPgjcw8FwfbDjAxjjrAYR+w2ha4d2g7nyR6EY4mQKa
FOodQacfd3ah6j8oC5gOujioxnIav8y3svzMNsiz+zIh2OqVoS3fcNNaaroju0ftbur5+qNODM8O
38iA4If2i1sYuSk0BnQS7mKJMaqL2oMJgt6Pm8vJawSF36eaG+svMB9oJ+eUJQnkqUMrCY3R2mQS
r3QvusUwPawldLif68nvx4ezxqX3eJ/wbKFNtMZONkL2c3p3DmuC332Jo7SP6ULDF17Z2JTo4WE7
S2HNwU1zEMmaxtLMnTkADZVT1nq15zmHNJGDPFmT6RGThI+DlgpCSXiwuXdaWlaC17pOSvsRQaav
JkY5VqCVpvCtnqZEwOSvALZRNOv0Nm6tsPfOmd5mpOHIITCvLJrSU6yff86znsiofUuDhr7HZ0mY
IsI4D0y55ag/YEtlZcg084Ef1RlEnWXD1mGyCZqzl/5xJNUr/YiUKx/B1G7R2UNAQFAK8ViZEFtK
hOvmfglq/GVIXKOdmyBzrJz2Ye/SDIBVqYXR7m11hdcECwB2oHknGg8NyLmE/ywDcIQ+LPDpP6IK
XfbgKjiTtQoUrmEEK8OBMwx+tjw/znrktR2yu1TUdHBsMDxk2h852wITmq78WLlMlNQCIpEfmb6o
9iEoJ2X1oaDAWFUwRn5O5BThs2RJTjtHBom2PsCpYOT3Jpx2d+ObeNZqAvsz9bw5Eawf2A5NThu7
o0mnGSvE8K4/jT4+vB+t1QAFpVLIuM2bbrlfCb357rrr8QNK4Rs1+NDMnEYsFbxlEs0feTNJJ2xI
WD5Ao0F8sJagjS3DCHlJig00YlA6CKTz/UezGgiOQ+Cc2pDhKaoJP3n7lJtbjNHAhPFIlE86SB87
l3aVUx1UGvy7U6IugR/fw5bAj4BxQsRGMHrlatOGywRH7och6QiZ5J5h+rBKmZzVB7U0wF6V5zRe
AI6/kK9e6oXHb3A8N2mZbnOUZqEO4pbdBcBC3rKlCF2+oR2Imms+qhoe4qTy/rOwSKgDIHAIIaap
zT5SV7C7i2rGwKBwSHPYXENKctz9aGCcggI9R6U7LJ94myRo3sfjQ60pN8+Ot5P1wdPohpSCgP7H
e1GcWah0PeWQcKy4h5aGSre3k8f+vBGryXsubaKezzlSimvtG+tmqhjUAbBU69shm7OKyF/UjmIt
pJ1Fu85HeFaxC+iXM3uLEnuj8r8qHX0gcYs9X3siIOizIM6eQvN2SfFEtOsByKOzFV7aVEcrtTOH
O98rOqNsNimdjyvlWC0cF9RjUDrMub7zklynoCF22DzDBwUy9PMwRTYosuTXfycki2HGbzl+UdiV
/ZhlBHdb9Mkhr7S5gTZbQse6cNVaXXB48sdu8rlPrM/rao1EHwvnwbFMlr+uyc5nDjlPIFuEkdDH
ONB7AnM/s7dUv0R6N3G6bQvMMnRiKaJIS1WVilK9lL8+OgmiYoLKZFDwIiQb3cx+5tvmt2nDPsJM
UCwnLBf7Mlb11Ci1MoW8cZAZ3qBHnw3sr76+Mg7rRvGdl4+kBbdKiTcwinLx6iNxxAGwhtMWSAC3
sBxrU9IlxII3b3i9d8MzNPLCh6WIwMD9PzZ5zahwM+8QCk9xddMDitQ0I+ZHqpTyfWdII6k3egjE
O25yASi2lNgq3+QYSKP8jylY7CV2lhZl3XhH2svRn03SRGkcdxMRoKJ0XlgZLJp7YqfWoFmxco9j
FX8+y0nXig6EJUOEHY68JgEGbpXGGl1DvQDfhrR7b0EFb0Ja5YkhN+ll8CSrUuuG7wsYIr946xs7
/JgIcLUqfF4nIBQGW+yKbv9dmZ4JjkhADF88XSq2+KRbR0jB/uJ9pnmC2a7minPGADEsc97iLz1q
8Iz3OioSx2NzTQSyaaGdYL8QbPyBMH3pmqDMDKUeeY5yAo5M1gbaBEB8vgErinF8a5KJ81yoEfti
S6wEBtLaqBF4cZw8h4LXi7JFBBtqXLrbXkFPKKLEuN+Xyl3ywfpGx3kGPa0N45dUhaUnneilKv49
V5pbeQb5oMQQ4QFq8VlEg+d+fNOBF1+LvECivWXp2I+hoPOSoSJxXyg0t6RNYfM2d1hHVgb8X4rx
fGUhvUqJzrLHDQ7b/iZ7M8uGe3Zhnt+xPg/v8uoqQWfPbbrH+TXynJhj62vk+Dyf4ORjkGoeAtBO
dscopf7yIHr6yallEIgKSYy563sY/3fiTGU48LJavLXuiQrJfUtXBUHNAVEc6mct8tLvwYwuY6Ce
nf+dVUDxBMcy9r2wPRNydU2q+H0cO4OxLEK87twg9vzgfRclFhuuVuU2LcQaDwAfNchIe5b54oDD
podf4s2QWv7w4jhft5uECYJRrUcoOBkErR0/3WeNDeV3gthW+tyDTV5/XhNURsYAMrRib8Pon0iC
V8N96o66Ig5QDxVj9sxb3is6rdRZup207CQK9Xd2wMiA2ZnBvSzinInNjfwRFNVoL99qT2C1K+eN
Og3mk+CErsPuMJS4FsCv1E4Zk/PR1XJAgEUZAGGXVyzWwlebGa2l7+ITni/EOSzoRkNTrtLZPZte
JLnhMuU3QaxxFVpZEm3vJ+qHTjDuSObniUUdGQb4EF1L3bIU6nJinOA6WSaNCXWhchIZlHfi23NT
kbyqig+Z0PWDlF97y9tb64H1toFX5sqNc0LIr4G1jAk336s/ZQ/7hcXU1Qm372lgcAXRTnVVHzNr
RULk7ZcG7lYMxcOc7gFgWe6XT/K1r+lm3LbhyakJoYLp4VmhLC+nns6b5/kEqE4F5n0Gj9OvokY/
COVdGIcJwHtkQlsEcwVnFYrPAO1yONQrna0YpZTH1m12XB1h7Y6N/Yf01KwBH1JNemxL9QifjVE+
vyYJRmPKP1IY42eYBQC/GHnCK2gEOVDGzXw4eKWMcq0nveswaUMwc5wlSNAscLmyYj8dyLZzMP3y
UEICnFPkCTwcktsCrkCEVkPPfOVPelRZdouuDJie0urQNTm9GKheQ+A872TyzqSGGWD7dd7NAEH4
XojIFajkSlo97wToaT77t98fMh3FAh+EdcMTCYio/gsl49lbjcauGbbTmSuERf9mtJERo7jPK1uL
BIkDhufpRJl1wx+YkOb/Q/473UT/KUqLuiyJm3jDk97B+RqiAPjKugRFFm9eyc8g7iTltGo+pEdK
2oq0dSyGSLTXIS/Gob+3gCWM2EiyclxBmD3RGeH6Eq2FU17HNEt+Yuk8M9+hwEqOuk9mSDFz15/S
nY9Ow0p7b/0Kn2SFWGtZ93UnbDTXBrw+zurHNJD6Z8bz0M3pNukeanQ8Nu4ODBcDhaaIrMwUMqQH
JpEuqQlabQUj3T3cyxyW6ABePf84ftJyNdpfo8X+2WdTC/Bdw/OVJdtbfa1IlrFj+fS93nICyW8v
eEC4wi1m9a43SsdWqX5QvopSFbc++DUUdueE3IRu+B8OMCX9jOxmYuDsjMLttn9K9xFMghb5y0fQ
wlawIh67YWLiLzcwYFIs4LfnKuZ4JQalOuVX0Nn7h9ompLa9qpX+YY28t/NaR0pYpSZi+wSpNdK8
1b8wE9TI18DapWc3yybnXgfY3HNxbheOWIPDN6zO6L+gtSsTUgIdwVeRkyIAvDiLtjjFhBfi++lt
tlUZ2f0i7x1XdJdHfxpjwHZVRJt/Wb3FF7e18RwAKeRBJ1dzjqUQxXTyz/WvVg1qRiouyF+FoWcp
RknOe6hTLU859ymLpajtvUClJDp3Vm28XWugxHykK8y9Hwzxrp31TzzmqAlN0++QikLadNki1k9l
6ztjX6Fs5j4oUsc/RcCHBwGWhpby77FADEnor6u0wloimtq9POTiBAk6In6JBS8hUffIRjpRFw17
DQDq6B6OOpFDiTHpVVPJlP6U8Px0Ctfq6KX4czFJoslnD2OgjN7F5OV8lzPxTNymvpfkj+F1XTnu
9PvwVlLAa5AN5xBEY9r1txsiWafpQJpSiOfX4CEste3k23tQK9BGFQ2eiMCNdxEVT5e6qKmAYhmg
XDKHkgwGeq8GLS4h7MovTtz5AIFMiNOU7ZU4L6NHXSAnCN2aMBsI7Scd8qSLLGYUtZyFyjtgekyJ
FmxyuvUL0vXDM8vIDxjRubn4YBaHqtPKL66k1J7lG8lKybQpIS2a60BMQEEQI9NgsJALxMaa3x9T
nIesvsw9LpHa+ZqNZ7QqT2fQfEa4C1zjwdvV/f24dEaCCSOHqlY544cCiPiAs0Vz/ENcBiD9CfhP
Cw8U63orSmgoJvXl4LeX+jNEhYvCaIAtyWWjGQmtzWJ/v4mpG+92sgmWFjbH8T2+cky7JB/jkN0y
/gL3A79M1VsXmyxc3HqQl0KR7m9sIx6I9IgfeNEhPquHAKiUczHbWQxHiNcvV9FI/97npO1BYpn7
8UZKIAY6TRtS+JqRK2c4a+DoAoXWYbWvFV/nyNAM1qfH36juFgbB7PD6yWf4Hj2no/3Qh9t3/Gy4
FmjnwotGh5/gLQTLVO2WurtrCvtxY4XA3Q9T1ISxi2rsIgEq2CMKOIXXi3mh/8rRm4IPIKfq5vIV
uTF+dtxLkEtszSwyYQ6KHdQgi8U0Dmu4WniYmLPfMY1hHEImXK1W1BNLGLKvAAIMKKjpFux9M1rY
9JulNqtsbJsrMSH6Tl2mz20gNxyw1y39x9WaVU/Erss7/tYxvjR9kVLnTPSexm6QccPDnI+t5UAD
wxZW8c14LdoB6+XA4s0Yr4pRI6k8zuAnwVtJBnRE+MNpDU3ZtbeLjhzD+PX20KG5YT0PGcpmVBdt
ESE2AI8eNSHSd8/vwQgL3EVP1J9fq60duqHqavirn+dStqZNTZRrC2SSlpyDvpEHV1zZ1Nr+GnD9
vWSKabSXzM/XIOHKKQDAd06RCU4HCgXrGQMrd+mx8oSqzgv+6XaZ/qL/VT6sc9/ShneHWQEov/TC
Of/RxSTcMeN/BykQFE3HCUaPmbHRL4hlMIKLAFQpOJyVXffWlFlnYgPqe0a6gPivLcJm8iPd60pk
SbeNEYZpbYSAGH5krzDO9sG9yvjepocm1qNANF44SNXvwo/RR9BiLec/SZR2QI6A4CWDojxgXqVj
tn+Fv3/r5C2vtp7tAn+2ZoFJiZZoOD8OmfQdCmZ6RhcPUbPJufTpz2kHa7icFXnqCW+sw8M1/4d9
r97aRrT0fTcYvLng1NwZ9PlUiBFwxfq47bFrt7NZVNWILFNC3L7/Jk/QMJiuT4KGJN/BXpKsYGMY
0N1Czt9Ex8mwQvkovsuvVrN6jJw7vFHX2F4fvUADUiIZ1M2hRuKXdF0ULTun61lviEp19gCE/uUt
x7M8iPLkR6Drcmse/WYRrAEu4aS/v9UMWJE8ic5WAKs/PhrSJq7W/pmDs/wANuhHWkPtVtvbqV5c
kYfz0wT6y1iAXSFTWGLH4mhKhTxNFS+ODaTegQ/OKlqAdT/oGFclgiD+PaPA0pp10xDAEIZEW52v
co5ua0mVYo0fiWsGnCEjj34WlgjxOOGwVyEedsFjrsHGXYyxrWK9i9MDf57sT9csemHIY/ObkvGD
mB3KjDPgIEbWCBTizRncF8KYMntLXpp4O8qGlFQP95EUpgYXw7Bew7fdvgWBbXAyh66pnDWo9vY8
yn5Mcl3voTpLk9GkzBYJzuuTNQR9WUM3as/sKJhgQ7qWf8bP/LzuAEJGbek29Gm06gyYnDJldITG
2z9ue2JQX6jmbsc34RdzzT4+lBi5DebmUZ4SyZSmEJhY5Ak6wB93gkNm8uaXQfS92aISokx23xxI
hTBOsciLoCAqnti7qFi1MCzaRRiwxLPJ2S1baUqkguaeUSjIYWq0uWJpTL/nJTqQ7/hc0aX8XUtw
cW5Lf92NHGOxyJ3g7J/kTI3FOy3n1fRWGOq4Nir0KMAdKLwXtS+GkesLcO6qREK2imKHrcmugxIZ
MFuQLafKdJxUQZHOGp54W9dXPa99DF3r9wZRYt5OR4EJz0aF0sr3VnmQNxalBd9HjyV8DkHbjuW5
G0s2YqzoB8q7CQlEvZqfLHg1viMashXi8gF9gjU9bD2FR6hvfULM8ZlLCEG2d5nmxcphlLMDJNJX
7flxAsL11EeoAdln7kJWEm9Y2ozYKh4EdCoBn2hFOTCZ9/WQvwvZ21JMTvtA+yiAr4O5gG7RA19X
nKJGJ/X2OLr7pPE0IeJNIVG0I1pORTT7iwo2uxLzAq0Pp48wZu16ePDxMhOb9meQeeMDFGLEWCaq
/8272gsAyJNWxG9VFB8f0vNcZPZuaOeSi18YSkGealTdAe3pLSNctMdA9Woql6Ln7akGUWuExXia
D95fT6wobemqPxpc8F9ter+3m2wjoYk/SEs3wqCl0VKpaEK9mgVsUdFi0RL7eCKIWwIE7foSAASY
rLd/3uMsUjw3h37mbrog7TrZ7KKYDpsaWE00vGTAYpOvunHqJ6/8btAag81WUk12+izDCy4RHScc
hwT6qfmVn5q+f0NLMgPgLp7EJ7m5I1/CLDNBl/+qLx67Ejh7NmOJ5iAzE1ejLREgm+9w0LoYdCqd
97E720XZch+IKRsxrFyXCMX7lVTOxhVv1WmG/kUJM/Y45RbduMJW/640i4Wo024Ba/0Tk2hUzlAs
RRrpAmez/hqW4Ha4Uh6uoPnorN5TNwu5whXZC0WZ8ky2nLIVZr2pb9ecoaxG2SLfIISUyk3GGM9e
WeEORNwGJQF7onpbDAZ24RNUXg8ZKqp7MUE/orn3v0rzKQ7773yPLL1HkQance9W5Gc3p4xyvipP
Ms1mzHIBouUb0z1UF1cxTszd0Mpk2adqPzWiC93so7Xuia+AatTHdKPyBJOLCkhSUiTtZeUGap4Y
Hb25dlsqCwCtCJvDYUMZHLbtfSq45Yo0emOVi6XNNbRuYy8sSj9zJOuCcB59n23VEbvrVHmIuTRi
KfOTd0rARWjA4zGE8xN66MqkLyoo56bkqPkNDwvlnhUJIa969dg6CFmWzNABAUV1bEpPxPHs641m
SwCYH4ePz2KQvtVbJSNbeR5LWQYioIlvVinHN9/RnnnGnesXymjtp7Kem6HIfR4PjB1/Z/Uma9kT
ql0sB81rngp7tKrHTwnybHyuBaFzLq+ew9N5jtky4iOErjfMfEX1Z6n4zgc+PT/a/atSAz/YTZAJ
7fGAKvIwlhER3mk+QrgMloiczyjJSXLRkydp2JbHVzZ8WFS2Be3iyufdzqP1D71mKSG9pYEA64LF
TnPBQAzgt3cirogoY9miaZHU8DLo3UL3fELmMKLV7QwI1EIqRpTNSauvNjSPrb9mRbGoXdyig0Y5
dMcNo4tqAP3dP6kqJJ5uE7f8UkmL3ReJmr77QAEtVp65vm032JhFc2gGjFUKoBwWqK2fGRKAjjms
619/xr3PX3NSzA/E4xrP056LC/JMig/u0jGH4NrWA/m5QEtWESeMC+PwLTddxJbFKNjSz9Fus7us
pR7Bt2Nj4mF6LFO/2SYERF0ZKzSSrS9kLx6yfgfJEI5cjmsSNATB+wPxlctZsQbNw1CXafSgoXOw
2cpYkuBJZlg5Fo2umildmFgoNuj72nUdsrJ9KTgDwtAUOKFzamYYT+JVDU/Rd3hRxywNnqdjlcr3
m184lpHx1Gb8gZklBQRaeW6g4jTPXQ3B2xOzrgfNOPp7/ZTYqvcOlC9EhiF/+Zg0swmgSMRBZymI
4rFK1GGeeIaLU8h3s6itzWaeHouf3EZXynzOQsTKWW6GtSa297lFH4D4xrSwP5I2W4+h4WBdP82c
UF6YJ9CXjcmJOZrG1GAfGgeWpxUA2Mq6EAz8qyB/fHJWUSES+y4RwIOZye4aOPO8yLJs0YCSRkv7
s2BSvjOZruf2Fz8w4Nvhb9l2TH1UO76YwL5aEZXvstWL5CgE0LqeXJHB8crDBMEsJzvny2eet4nD
kTm6tbjDmiWlTd25Kvbl3im9hCTv8bFNZgzxv+2xFyKB/6FZVe4WpkzMCwcmPA4juYGEZ2o+xifS
XB9TpUMOl4Xy4cwf9qeGz86nx2AP0pbHkfrg1xXICUGLdQl1Hf5eRFvg4pjReGmTztB47EjHoaEe
GjMDP2wAX57xxiLyMb8G3nRNgjHMa65L3Vp9qkYfRTay9P+ZoP8gRt1caa9rGjVRbgG/u6Woz5Rn
c/IY9rczji1gpMRIZ3FnGa7ITAPK0tJSf7g7V1JFMKj7DPo26CgZvkRIuN4hwLAGu/p6wEmvcpTQ
pZEW74NmXeE3hRfNfFxAMOzD069WSkz5q/xsQsMs+J+4Bp+sYlE4pTbYsfgSivoev9OGUeSJqMDd
tnlsHRYcKnB0xLsLhZgCtKEvCTxFC6VGIjoZo8bwTXIKl0xxv2gEfHtpewBLMDd5FijYXDO8pGkS
f59Yk3+l5k9UNY44RDiLVE9Hc3P7qTtJG5XkIp95tiGsDgXJcfgODjlfikdNjiJrO5D6ni169NCi
iedTHy3of58MPb6jv6BCP28hJDk3NJFKDemRwftUf6SpiXlh1sNAJfZlh0PvNq/fc8OJKSH0nrUx
0xtAXpg0/0Jpi2aLC2P+qyHy0AtG6Gu+/blej7nBnY+9W1MQo/Atp0IwHBB3uYpq3BsT4ylPoeCr
gUTPGkYCvP3d0ZRA3RzNznso86DAjw+An0T34kOpdZ7DqFLE8ef0iVU9q0SYjGgn9VXJKNpAqed1
KFHTB/a98Ll1TA7J9gsvGlFqbH5Ab7ii5n1XdMLtBnhqf7YSkfyTsgF8qgNhej/WOuwxXPyUOMHX
oX/foGUaC9UTyt32rRvjXoK3Kid6pZnz3eayxauH6kH5kvksQwmKKbsaI6ABJseQPhfycGfeCK1m
vuiS15l6Nw1wl7iSjxFfapG3OTdkaIAtEUJ6QF5eLWe5gwi9QCgLxzDobh4EUnV/UsZvcMEnEwJE
9t7Fdn3M450rIB2BG5TTyGlV+EmTEHx6UAKd5L/59No8dcgAurQztkA8FjGTLD6Z6ROdrUjeLrzP
hh0OBLOAr1wMypN95Rhije7NjlVTne/V0sHR2Tp3YCcAFIeWD4j6lZJ3hZOSwhPs20+Iea4/Glwo
sprCdcDsdik2Foj6sNBTEkA+AAglgh54w+r84f7qTF2qQfMwe9+oMcPMkVEGS2y1Y6BbOgGmgh2t
1GD+vmoX2xR50pcQQ7oo5CwVevjFONNpJhk3N51sve20Pf/e70PPd+dZk7m5nKFzB5k6UKOgOZ0/
fD2e4DPMVPpnRgwEpxbyoTxDG2fiTpC6ySMbhMIPyv7KmWRDQBW1F5Y83UEc6Gqg22p+tqInj26b
TqcFbMnyTTnV7d+ohQwRqWrBCD9m1/8zqyh26ntOIazXhjiaKe2703hgwkSIWRahptwlwgM2CAeD
BAP2xGS5K8+GwY3c1Hr2dvh9Ore9t7fkoSwWaR9xHnfuQfFRKM4pedhRQMoOfPYYtIbUYZRltJpB
MC9BkYPLx6qPi9pamUITYm2yk6jBbUIGLPiUc5Qc69qWFEGwp4DWy0A8GLZkGgLE5DXn69rxFJH7
3BE1t3o+7YfSCaHqQoxfisKUQVvhotz8KTCfRcPoN3Q8EE960jpmK0t3ZpgAFsfGwithUX1wZb3U
kXBVI8cazZH3n8F71kqN5Q9Xl02SbagcQ8y2A6XC4tbU72Gd+en3rByycLcO1piFrJ26H/mkAZzl
vRClN6FZargCgasTb/dDOqtus+hC+T9xqRYlFmWa/BXbBLtMfrRbLush6sXQboOa3tqjSfqNxSXQ
09RDj5McGfKDV04xx/sKfNrWiOsYZUQRYR1QKdmo1iSQRWgLHwwSalDxc3f5I4hUxboDwMaYa1cB
LyUeM5u2I4lkoKbGZpo69oaylDdnq43+wW9TUGEu+ayi+EXOX+EpRPuP09MJKvoaEOBF8/Q5YHgi
/EeOHDymC0pBvmngzj3a3V/m461JVuPVB+jdSiESkfIU2gfk4hmD+z97YZYgayI10/uZmFcPLDNt
u1k0wCGSQMbmXwDrE4Tyf3mvswOsnJ58/KuCZ+R3DLrWCSe7LShyVOJsfgct1oEVcJMKHtAD3TV7
jRH5QPTU+3FW99xZc+he2EkwSy4ZMLm9HlOL/9GPTHkaxb9n/Labsy0TirxTurh3FdcbvygrB7SE
tQGff/XqlLYYdgdBEqPmiSdSOz61yk71kicob7yRQFWXFFurqQXEX9gYzWJn4BnRWLu2LcKlQFSg
BMgf2LdnRkcu8gbpz6vnEeRaev4oYIaDvndj7wMrxLD6t/qgq7K3xSAdWrc/LuJBXKPW8jB2anqC
SC6qye7ubuCq99ovT/AuzB3anVVDryQ9raIb2+E7Tcx1tFSCxaoQ030WvuIZS8u5PsaKXAV1e8d7
4u/rAkc7JW31sFBFrP0aXHSWaGi5x61q6tstl7Re2VBhVEfoMCUf4NKsn89Gs4MQON27SbxpdQ9K
h9dICiRfJ0NykbY9c9iflaDoDtgBCSvmGVgnQBonuF+ArDY/aoOPxW/vTTadCDwY/Cs3QbL9NErG
M+o/rRisGmpNZaQbRjwjp0TAqeGyZ30HCOgGNkkuqDAzJIUR3HAodImvQpNwO+Y5okJ2yzw12K1Q
vyFCyDfKSAkpODTCxvhfHuCRQ/qAxB7oHWAveJDXf5GUevBBDVwpa7Z9yWvy3Cb112HJdTt5cXhc
PbGtUoOR/86KqD5pDZMG1Qhb4rsX27+Q8c1vfv6BrQxOr95hG3lMliWdivkVXzy7GtRp8EbxQNVq
gYpKziT/mfBT/kv7AsdMJ5zE2iVvnMhxRdzjHyF8nJl06r22d4KylguWG/EBE9GI5B6VIpesiHfh
II4ewAkeF4S6KLvjqqREUWG4CVJlxl258jLd/2pdthq/YFVJVtxfDUe8lSbfHJr2lIJUL6OM4fbW
6Ilh9AX+ANJIADxiFQs9y3rVGlf9Hk5ZxlTvpwH2scs3zi5xXb9TnnDsKj1RAqWcLsHOsh4q3kUD
pxLY6mib24+zttmcPZXQ962+6jLOAyzi6ZOSX0ve0wF+M7u1qRPFlR7U9gaKwwi5K4Doq0J5ELVw
qm4k7F0s9YEscT66rl7cFqKGNeEhg5RfAV+renKlDTSWG7iOOU1ivlnW5E+4x/PQNUbeQrddhnqO
J649DRpifiTPGgCOgRG4Cx4BYYF8HvqAfPJ0H6dxi/2LbUclqWc3Kyihuq2+4LHe1YxHmmC8sb42
mWgiBCKOQSP/v2kJcQxIFxJEjuFE1am0Zz2WCTCp7iaJzlSi70qeOjk/tlACeHbWBOwwBR+eGvYz
qmY1roFmfmBACig4U6pyYm0lMGIeGpJd7/j+s+rE1/XOxcfv4KjZRboU8I0OvEvz6lEbra6P6fOh
JCWV8m1yI0D8duI7NWGr4Wv7H8o1c5R+SMYgpo3PQnKYU3rLc2wYtXss/AgdRuIAxsWb9qn9aQbN
CXjh8gtTDq0iFXQMDyHRyR+3Lmle+sT9qgyEzuNzyfAQ7/n2dTUhJrCcKzVy5vBYOwPKB3FlK1nq
jkYFXyMvNrhNFh8lGuNJYMj0dOKVqNqq2u3wa7XxxoQ5YrykuussSPEAgfQctbA9AutbtJ5Vvv7W
+Q1vSkIUdAHVKzAeSt+RhPPPrINebNok+NvL+TXwpU0B99y2jBJqiBs/sxJX2upxPG4s05UOy+of
kkcgkOT8UmWZpEi3oWIc0RPRbQEsmI/yU6c2CoCHo1kD3rdlhSOK1QuRLbIdpL6Dn+rlwJaclcBH
uuCNLr7bxyTuV6vBAeAP2umDlHnRhdz5iupKkz4DHGcjPlvZBYPBksKjARDCqBSs/p2nzeZqoQHq
WhjQsubpdIsQRO4Em9GAcM2KcLwOSA75Aa90Qb8PMRDsfHmtvm6OBIaef3qxrwBEJDIOhSwbzWI1
3O+vUxl+15F6jbURp5O8T8VIOj1OB5orTQ2z0/uewxXrRPGm868TlILIDfAtFGwho4b6IQ0VzRav
0G5yy3sWUnskZ6Z8mIJephlEPVH5Oqf1RXLozffHLHpx77JqknrbqnT+QxHOeHKxc+UxokdSn1ox
JiTtjK2zrzswIckN2zFyZyNBL3WemmVF8r0A9s6ByCbsH8BJs+VubVFmyCPaDOmq5lgUO/o8Cfss
vpq6qoY3VtaQA/v2l4+t/zvsLXQMlUs9GjSgzFV9jdwczqHUyXtEUlLwMDW9uIsOePCrJ/aGnBH4
fpBDAPdvWO5aUwx3wTQJYjl1kXrQGQypexGXBoZItEHeMgPX4RonLimUcciFx7DDQ51ACeNu9+Bb
yEJpm6VTYGqpGb6ooGoavHX7m5mVxep89maJFLIyfV9L71g81Iz7J+LX+TegmuxmHOqjbBvrkwaR
EaUZkpjUrpCIGe1p24ZC50+fpGMQaZwKfAjrwQ2joxO8y430XVxiIIbnG0B34PXRdbV28AUj4oM9
HAU3Fb/aiE1OC4THzeTnN46sknMjIDwMNf69p1BV01JNpBWY28f8wyDFx4/SWuN/g3AYHonLfmH4
esJbmD9+JLCt1sEG66bBQwPa3e0UemaMKr9nBkxibn/HtsW+dZkruSkn/KDjZ5iLOPVT7YZ4Wr6Z
L2hiTudefQQib+S28YGxadf3BFClA1A0YENNR98dzUqk67WtDtto1tGsf1HGMdgCp5joC/NDmGbt
bPqeXSOyteB1wYoSRAEBZc+AlMlNIdQYrBcR7SGyV8ne/o8JlVS+OMMmOzPTS/NDn8hFmd6Bz1H/
O2z9lrV0KVaWAigiviZyUhYAEFkRegewn+KJenYmmLnlpT+6Wpbeq2mqNvo+qH06uvBNc2y7nIXU
bb21+tboRrHzbAf82MYYorKNdUTygPk2pwKctO8uxUw9j+CeyEDYA/Uk4EhczSzKRTIRcJcuolT6
pHAQFUoP9rYbb0LwerqHvGJC6TDE+LFae1i2hkPCHbqLFZ8yXYEMLrPq16DJ+FGrY2kEgEcpmV1v
I5TsKj9whcDn2BTMmyXMlgra+aLzGD/sxawNztUqUxlq4A/85Ijbt5pBA+pBYOSRluO14IEVlsA6
LpHIb7lZ6LWynoadB2h6WmH6Bi0geuEkF4ouiIcJCowykzPZRmw7WviMYzzeMGN/0pSIqeTptk/2
yx+51iuBCNbz/2F/itfF+tfM7YVi/kfTy053nKM7Gum0qnZURVyzP0qSNmId5k1PisBO2zO2sx3O
Ll+bQoV8ZF0xclrZusx825EJ0ixjYwvbJ1DtulmwJxdacVBQ1qDMtPt/bnzAoQht3RyCfpRjr+ue
Vd0I13orrjmHAahKEH3Y/lFt7Tu3TFvQROKwqODDxHSaqlAJdlGtwtDGHgyje2n2/SZ1Att63RS7
EPD5+UPRYilKiJrQiH0C3vaX8vf5XANkSnfBFvcIfAptMcoDx5v6+h38da23cmXAivX0ViiUt5Iz
t7JuYONWoItZK5fgvbiQc0t4663InFEcBRd2QEuPJ2pnHQOwBpf5EnTLBmCvf+Cs6wVySi4xI52b
ic+eSyyxPPGHxu7LCIxZ1ngyGVkfmXh4GaCfv0XlT9sn/SNWnjUwUiWMEwRZoe6wi/ChvH9EKnHf
4BbopEFPfGANXC6BuTwvF4VxY9RDDoyOAFmxkn8S9fScFpMWnvTA0MFHw+DAIkBIiAh8i1XQb8bl
TwLCju+ZCiFqgQV9l9e8wcBiTEjcfscY8mRFvSTheANjq7nO3vqgpFwDmdv994IrcpVNl+U/WXxw
Z6ap6s30egJniUGJzy4lvOLNcfYY/nulj3Su6VhNDywOHdYw0owgyQofbLg5ryxHVDW2vEeK5N72
ENWoF079zyHU8r0qnyi8GFKbmZ0q9edRrfTrq97G3ieKAomsZmK8MuWAOtoBMHpVULW+6JV30ZdD
WJas/VV9nnbgRp7W7XlgSv7qdLxLpiD2UwnHZmNfqMgejMcsZ1OABIOjZoAXDfij73KELpwSBa2s
REQUeryDW31Cm4oeC36jX8jnAz+2chnh2a1bhoTdAATssRGdgGv8Hdlphi56eQQnpJBCSSFwclHr
sBl8V3V4QRt4wEwqAU9J+269mSD/+ZG1gCSQUtJdyuCON55P1BXDA240iT6iCc56bPAI9+65Sd7q
BFNsEaMqKqVpDYK3R3Nq5XAcNdmZIjStdc9uSclESQ4f7x/JOdd1ss5TfBvG2FIvo+uwEgxrxiLk
p9O43NzhIKr0FZ0vbX7/fl0KHMrIFW+bSAU3ZPNm4mj0ZNiThWT9O0rcQ1X30SCVJHMORJQGZHXQ
OernkCRLVP47FFSKYWzar6svIJWa9LeqQzvwtQNWF9T5PZPqy0+8+7Eu5IlM2f0pkKofvoityu8b
mMhykPFqe2qIvaAHfVAXhxlfE9XUy/xKEBSKQnIQtjemE7RchW0UrXwbKZnuntF+T710KEHnz4ty
xgjgunRA0j/eWpkJlz9Ra29dOyh03CqiuhUMny8cNOYBqjF10qPXI3bjxunv77KIpSy7HTzzdPMM
vrp/jaFAsYmeeYd8gWNIREAvPGl4si53+Zv1Tpxrq9NBM32v4X8jdj+QfOD+uychCN7VAYwJ/+T8
3cs45y+D9DCwFkDJRqyCZiSOcXE9O5AZZgneAihs5V5tNpDMjELuU9ITkEJfdvIBGpLRGIxRcyQp
q+VOazJvWex/l2Id2pMwccmXSiCVPZ/U7QZJnqg5OKZKbja57JIWLaOueCt6hO+iVYzCmA0R+2nK
2ModVA4L/eTc813nOO8/z/26CeMKqS5Ubmp8GJL9X/l7AT/SAvNk9EBRinVyvdJKnXOTBrEBbbpH
1JJM7ggoQ4C2oi6QcUmOurggV/5NtYLVQ6FLKDEXa+lHgoDFBBZXf7C1t14rK/ilQ721UTbOAQfJ
1XDy/HANr2kVBIUSJ2anvhhXftc0eccZmbuqvHbd6gv8EnbXDTvC1BObfIU4708hq8CkTnr7D4yP
sONgXR5g1pnGiwk4SYfb2XJuJSi/TB382cz7ar3qUIeJcdCB8b8ml1UMRDg4sIfQB8B45ICeFFmz
q66YDDXk1mFImrQbq0wZ6hh8u9FKb0/nEewdKNC2GYMvBnTMtxzruFC9u8YvsDNL9wpbAe61w94Q
o2TYfKO5UXQWxgyGdIE2vny3FuS7Nla4aHj83jH4Igrlz+96jYxlvBfwc3xLq1fVzv3nW60C6CFD
kqOUJ/BpEI6pDdbw/sxOw7hnESCwD4P1xFUqJ1H3xP2FjwuyhdVCEF5MrmYQ79I1HtpyDHxmRsf+
jWboGAQXi18rpbsHvGivVALezQ1A1cToTOEbrW3bL06+OumcnxopawwcYDWyx87haf2Wo7daPqNR
aU8B3X/+MLpqN+fcSZZ/fR5jB7liW9gC/ikbZJe6X270eWP3l+Tbt+IJ/3+F+oCMcmZ2b5MmyvIF
kc6GqnnXlBgSjHvmVE/0bBMgkI/bnURandbLApjWDQP+N3/lQoTRmNcsJn3o37cRM3HbjHagFnfA
/ptpThnNvHHx47RmapxoLS9em1e0r9ZdwH65mmaX1wajDSu3P1/UsdWxnIerYmK3IllfLpwwdlWf
icvy3dn+gbh6jGfJZt6YHps1txCbRI810yAg7eqKcCPYOSu1TYbU+ISy4qSm9xgGOJKpfwVmoRB9
LfNrXb2DKx3p18uyHc94VdCKRPZrxg7CG15wLRXUdNWGKn4fmMB9lBPvUci4HQReLEKizvWLW31B
CTOZl5RZi+pGNwEeEA+RY76E4o8Qrbh9qP8/z0oesEMKe1gwOl5sjMAtq3A9eDTGEaBHGlAbZqZY
AqKXeJFWFGaKwHJkeN7qe/pf28HhoGWLAkyqDRfglNmd2rAvlw8vDFrPPAAgySOXzSsG6DmD84EN
jQTHN2CLNIyQ0I7G4Nddo2L/MCHC/eTHAL4mwNcuTF3G5BJ/o5/uuPEp5Jg9QbDBdN/R58ZLOV0C
+vbXOIG2ieONvsFhLm/UBwImA1cFBtG0a46ajF7DTzy97SKE89hqF1Bht4swylzI4WHwAnO+3o3U
wibEyDFvT8MfotfKAkAqqDBi2R3I9orN7llitYcGLI+30vVgaH0IqJWLmdBHb/n9kh4iLXNj4hML
x8jDvDwiokLChsBrYXIaGMeohtUErS2tM+UTwRWG4SS1KmABHqwl7QaV54xEta3G24oonnM0MYT9
Geezm3obXQv+LvbCkKdyE4jgEA94TUxcMy9mJzbLhP+uP3bg/3SIc98aVUJVc8IFQzy7KAfSzrVo
LiOQoFj8RNWN9g1ZYVTokqO6N5CFlG0r9g9mej2ZMz20vWRQHfJMBJZD3+2347RFv8BHg5imL8UA
Glex/UclijjKwkWNC5k9TKdq9KpKOTgvxtFidtPZ9uX14Wc7orw7yyH/wp9spLnsv+pihw1XHYyI
ZZ0900WUBAnOO74w81HEAALuOvrKDq9Bmpo9rS2LP8XbTADuD+jgUrZIpJ4pDmolUl9UrtsOwcOk
09+R/VAuAGtB2BRJQvuwohzUNW07BBuEuhNahq5iMPmZ8XCo0v0MFlsVhMsYfJov6RNfw0ABYnKy
s5cEkUv/zxqZNT6MjpzNk6oVy7O5jQ+ymlps03Qb395kYy6m8xiQe4C+ugMB2+Qyk7KZtHJ1qiWt
M0+I0AddPR6qjg1fGH151nyJj7JfddxpMfFbiCPvFZ7xto0DBOKgQETQF85oAad6kUPtYVDlKPST
2UfuThb7oTte7P2REgkcEuUQ75/E8h4FmbFf1yeKLaOMJ7miCA0mEn/wsw+xSMSjYvT6642+cUqp
DHopD3khWoQLqH0mMxe1Ub9QE/5Oo6Dg1M4kJNrtbsIIjZ69lPROFk9ABi/5VKuQ+REFCXZYLGrL
X8x0LMMX2fkpKl7AUGjETSfYE12V1ckSSr5tQaOZIdANze+s+MYRlCLjb3ptyQQea+Zi1SimBQpT
xJVjQ6k9DQjIqmjVYE1nz2fo1eSrpdERdvh8E+IuHSA7nEMZEvWQuB42j9hhDyN3rcmfVIuzC+Sa
awqpMaNbUISdEvrskUe2VteKTJHYPcqCCl4k1J7AaMviJHNPp7VU/FqtohAN5a7A43x7Rk4plNDJ
SiWKTo5ivjjMN4X7NqjWe2tV9mJZLszZGTFZ4stcW93oGxe7qUwrh2plhmgu6mOLNYKs6Jg5LHHf
0WP9lhYQIYM8UCJAADajNjqsZhDSb0k5/qXQ/16ZlP0hf1mmwFnFVOFszNz9N3IQcccL3u0EUSto
tmvzKu/VQQtPhV/UyP9CIKJiAOW/O6tNDPwFg4JNrhd3bVDVUGrHfwDiIDSAz3lVOzzZTiqgO7Xh
hv68TZWnGyYNlae4KVq8+FL54iRBV/Ldi7EGMeG1G+gK0HliyZm9XTp7phaF5WmFlxtWk8Rm8y+p
jy4F7Gngh4ZFYkqY3WY7lWs6k3SUVtGtvc5Tf3JDlXpzP2DtsiKZjFBa8QruWJd04WzeAN6b0nHG
YB2GuLIv5TpDb7+MfQ4fS5fDQKYXdq/26q9723rCYnByLEqaWpbIsjL3bi8jUrNZjCZjLoUt5KHL
1D+11mbznsWLMcbczqX1XpXdu6fVWBsJtNbGoU/hufc7ZuMFvq0mRfItCyJMY5C2AMxSmUm+YlPI
wsaGIKSyebWwBbvSBf9XM1OuquRscfv8AE9K0cWAqmXVkq4jpQC0kHgVExtaAZIraiJNSnQufHMa
ZSR6Efgmr7mvh2OS3DUoWQBsfmk9+K8GLpZAOSR9fllKY+jrog3yKEipYBsXGue2UWBi91nprrs4
KXAjFeI4Fwtsd0EyveBhh0cixRBT5D9a1Ss3V1B2Ikj9VzMl161v6gRSnuvTcel8/Q7zNOX30D0C
pEZPquhX1Xn19kp37RJZPBzD4qveY9AEEZoGF/vFkbFAL3PTKsgzjR4p4o73r5TWteZnmwDYNAU4
CXL6xTNwMq6bT1yiDJhBPZgVeTBqzJlFHn3oa9c1qL1OzfkIPTesWVjh8jaRdiw/2OmFZHi5LQE9
Dh6F/PNfNWXkdDE+GN6romh5yG3iePnXt4vuNkGfKEEr0j3FUtvofroPWsZVGAdztGbKkon6XJMv
pNNVnEA9Rwj+4Zyq+ZdSroC1pJ33FggeqAGatqEenE1dOBS8+GUDx0kQPX1rB/I9kWvp2TpGILYh
CuED6P1DyHswqrizCe6eD4kKpduCh16StlCPtJaXVKB4H72XftqRfZ0Zfvbt1PUvo/MpCiwJQFuK
Xe0D5/UFKM55bAyNSijxXKG8GXpve5gI/2IxNzoBwnFSvqAtWciMKEmJpbIxKvQA3wy7wWUXs/jJ
o2H0mBMClSbsP+00NQ7pWr6tqsrXtREY2sqpDAAp7H5k7q5csmEY++/6IFzZ7r0KnJOAWPAMmmW0
Hb2HR8K+p1jtIXZ3OPurFFs8qmbPh2opYKbfFjksJldE/lpsorjk1/z2D2EcGjkG4GloHj9CPiH5
8rJ8e5Jz5U4hJg9kYDgdE09/R+oPpbzEzL9HqlSdraEDjlBthbJK2Bo3KW+vxCP3FU0uOig/uWY7
p2I4D0T3lWwQ7s6rf445+9Ut+D+WAall+EkCCjh3optY9xmXu7XiC1Bix43MsJB+KsNaqm1u+2y1
QECZVknGtIXIeNmcaMyWyIB68JeLXphl7VJx3Fs/jLKWXhbEsz1om/XE6DA/HyJ4f5lTzh0Y44BJ
XYl11T43qsLe5bwPzQCUfeKxxWrtn0WIoQhlNCM9ZL6/LDdsVZqaV/ZosZWER7oe0QYqiOB7EgCE
WYiaon2dqYHLESdJFP+MqnYnANkHBNQ4xjcqB4+RnNiB1GdgAkp0qXH8z0kYUxrz11lerYfFVj1O
nKgqRaxjBOmYohUntZpV/8hSG9gCjs6n5GQ15ssR6QtyWgtyTCeKqIz5SufIT2E/NH0ORC6yL1bR
4vNERjXkXhaldq447TRTK4tx3J1+JCB2hTj1Iwu6YiqEHaFoqqn87oMVlDuacSXKIuo88aAXjDCO
7kec86AYW9/NJr7GiIZF2HxnthqU4hiy55/3nlndwP/Lj4a4fKIIB59icVs5K3fwjTVQX+R7YDXS
eDeQqtB/4khywTKCadSUGIv/gqQC6kgLp6Wu/Rw2k9rbwhUCH/Fx65EfPhNiPkUO6SGGA1wpTYXe
3PZja3Ad0NHPxi/8DB/f+aFQCuh1HpadUoiXEjs4taIng+Xc0C3f85BMXR2wLWdsb50LSWeBMNd7
luSyLhqvaKvOyOpyiPIsRUhcPGfBBPhA8B+E66jkxgPlYKxJ2KVnKGeqpXlfBTVZoo+Koppw2rGO
Z5D78Ex3LsSoX6t8yS8Wm5yeV+R9q5vIX/aNDFxK3jkrA61dLRB/zeG+s0oD+AGOPIpoIumvQufV
gWNVzFRkeq/NG5NyRwD5RCy9rjPRbhK/T45NrM3XQwtBo19x18GYSq8X5mdPP9CwvsxscfRfbvhU
N2gtV7iUCSi6kaA2lSrRMASHV2xuq9zM9cPNxwgiZfmQzdOx48gkcYlLkiHCiu4wXUxbe4XVJk1T
SGXq/jLlLwY6SSwFmE9hf3UCBK0Kw9HRe67GKNUlVQhmutv5/L06wVS5V2F4nO28KR0T2duo+ya0
VodQgdMT3rsiPM+lL9ujkFl0pHVFQJ5Y6p8DJTMES7W7g3KcM3XVoSbI2VVTnbDrRfe57LC2ItP6
7I1hPeeUr9SKPNaGU8pvTu0OUd6lx7Rj+EVYhtxyL4m42hfWemt2sVLAQoUP/qwI6EVocl2wakFB
ImothfLgg7DbQX3Q53leQ7T/qtXwek/hFYs8f3CCJcFnyof/EzQhvguPEcNdREQu3JSOqVFKTClB
AWXYduyHxE5lgyAVIqayOanKv0Mgi8k1scOA2v0J4OnRa8svebZ6bkBpr+k/xS7Z2V2ZgFXp+w9i
NKzU22DrT9VnplN3zrWHtfHdZooMhNQ67/gdqRG4iTw+cnsJnTme+bFOCasmNhgtlz17jSfuXsmr
LRpH0RXj3k29eztdlAO4fdjGVD162cg4IF0hhzyoWh6QHWeeaLbuOgHHt2bYmq8Ec+M640SVrd+i
PtgnQGQ7eW4eAWV3qKen2i9rgzWuYeqfodrSkayJlPqbDpAxyfOIx2J5ncUB2oo7VaqC717Cf8cH
uUX3c2KsaC8w2hlgzHjBGkB859UIfYv/GIiZQrc+R+vYUskSbkVmM5VMNU/aF46T6p/WBEuUauGA
4ldJo6E6OYB0lfwHXvxrwJAg0F+3/0r8ys491TBassk7c5gyDbhyYvaEZFeWHqWUfOQN4TXMja/D
GaNAZ6d8YvdGgmer2aHJZjk4VQ0NVOJPa46WiwS1U02aVjfdSxflbcVwN3K55sKf7qf/ALim4fW1
GRNEOrr/Eos6ZbOBO/91K//Rec4UJlpAdYi4z6FdxB0DqfWLFWdlMB42lMgBmJz4CqRbq6CXy1xc
5FDukp+RWiTV2Jg5EfM9GS1vwFsK14c+GiYfjZNY9EdFN2zVcHBusqYyJJnWX8Mr4p8sxWNHNa8I
A2Aq7nCmjyionrLPJEkhUo/Yb4mGQC1A7PF2hyTdwswhH0HGylA9Kuo1cDnrdlXRrJ073DgDljfW
EiuPO0FEL0wZskQVdU/UemhFcLNqG0GvTITyLg3aiI4JbqpQOYvmvxFjN/0YV3mbs4cnA2Sy8zN/
yyPoURCQkP6i7wT92IcaZG/978vD5qiDn7313dvnFEpDqAKq5jmbWWB106sEl5ALfBV60wHaXw1N
nRwkrqLjVIdemmqZOgk/3qjnvn012+h46V3U0tmqptXCLNqGvHuQufcDmC/i/vd2KztGrBQDonsO
OM0QWn4znhEX9yDKhmZCjrQS94RnhEdHWGF0OfDhB8odNTH5hxo8MbaXvD1Ikd99Q+92gxmbXDS/
fhhoW9yGSeyThjflRpynYZSBq/9qVBmfXHS47uKrW/ttNanvaVCh8tLGZLjQEJeYTWGO2JSaM8bT
ypykGYp2Dw5RAhfynRh1YLi1xxMo+7RokrcyjssIvk5l+6PjeX6+CL1rLLBG12IJIWKU+AST3Qwg
mS4BlpqZGIU5M8Dk1fTdvxU1028TJGxC62YmrVUZnpe+ZVP9TXd1iK6udiu0zqKLdB2UbJZjYh93
AcpHg5dTzBqY+2d6yyzNlt6mzy4KdIT2xayMaHQ01STw7IkbmYyr3aovak2NVUQG+SR4fB+ZvOHT
BZrCc1fxvZ3DUKOHknOCbx/I1KlHxIlFeWNTKfd0zZYCvd1xqtTkRQIL0Sbf1hR9MPoYmo/7gD9A
iYOyJzxwt3dv0QHfmcNPlIszG1FdCzc78gjkz546Z3ZXlStrRAutxbUNWhtyUKnHrskSBE6bprCG
LR34fzm6OM9+P76R86wz9pNns3TjdxazvVluhVGb3hWE3ZpujzYdThGSUDT34WZNhrjteZ/h3YSE
SesCHHuoTDpZX9wSSr2nkFXNqyXVoLQUou5V6U5CuNf8rLMgubSICQiRtCYU0otFWN1fvN1ziEqZ
RNJVcmsVHb6jweUuFksjN7HEqNFJIOjPK1qA04e+7aKhUHnwmJCScv0Kk1VhTwDu2gyoEufNqrRM
eBOApfBgNs7epXdC0EUKrbZLYxZ77MrPBWip2gBVfdZQv9CO1Xd8hGNAw090vCFDJtJyHm/1FYvb
QS8u5rTUlOzvj+0SxuGR0chg2iAvwWA4QhxL5oeBjpo0n8Z0yi/leP1l6Z9Csko7vOD25wCPD2ys
rAqNKKzV+K8Oa2umYDcqDw2Z+pj+Oxl3EbPhrybfC59TWEjgQkgUvT4e0F2/H4tJDysGZyl46puH
+N+3L67l2Bu9IOOta2AxnX9JDBFM1o6qgNan/+hbtJXd3vydfGa0XFe1cmlTqYbZ8qD5vjnLAdUG
DFRBRV2g8X93XXexR5tARFbiRTDrzsT7kezEoyCTBTKnlbuc5BJnpcHNL9RyyCz/gY7RlPfKB1UY
/rt3pqCtC9KdFcWxHzBqe5smKgwvdTYNUnttl8y2eFlr8kBdWdz+ttbwh5/t2PrbDRGU/52Uf9rS
hLEXxSHQyB7LWw9YTbvi0MQ9SwC1wodR41zutwn7m3LTDfi3wLnm3OTb8yTw/DYxE6UsZC0wsXm/
gMhM22NTT0xGYsWGMdNS1DzW2mJQeSdZg5XTuEVNg/TM4rDHrd48mDZ7Ik8z+jVPswcMPyNBPBMi
bUhtqAplmsyCMrpNp8d4MeI/AXX+jxB6r12tjEKa9zWixm4DBe8p7rEZOPFB680wHQ2H1upSFAnK
6me1lzMbGKbCDOghye79Gymeb8G14iU1adXVedWx8YZWENrxCRnCy+4SPgd91jUwie4aVd2Ay8go
dkdK4gYEgSMPqQc1Au4bazpXHWbXMHG3qr8YSIf+2ffIpwzMZaTtfm/UM57aFpecAUTNJFawCPbj
4QpwhvcH1gI6Vg+wFmtqwTW5usJG9Up0BxDXs/IPcJWuhoyPE+92SuFqRl0kPpmORwu+CDk4mYmH
JJMs1EiK40+DQyyRNu5b2I/cRv3DdNu6kVAilOvnwkLdm+7o9d43ywFgV5kLQAM9XpN5TMZ5+Rvd
pI8rSPbLJvXO6HyFKwcTBkEvWpz0+hYjvGPLEW3coZSnc93bpGfhCcKApZ4gnPLjcpfk32sWw5OA
1c84DvzDOtijOOVDnu1IMOXjpHihUaWEeuUDKt/rJedO2nyI0mxXNAbe9B51/M1IrfY9d9DoWiPU
YFtkK0JKlx4y2fgDPCMkCJ7byJr7ikwPVSt36nn93PWPZfKPYAqQOSp7w/LJH210gdCCIhH6TtfU
gWb9gcGun6S8bOlp9RisMxXKwD5socUiftpGX3yFs3hjGvthUqBu+78Fe084rWCY3o+7flWXOL81
gcpo4GpGIuIBDdB86HvECFs+DpUWiSNZpKw8CfD0Ql0m/qdv7Yws7/HXsRshIz5hvl9bwDxXI6mA
MCZiJmIY63ETYCmi12M1P6le4Sx/h2FkXe35JlnNOywLFywQQad3j1hYSP5Kprt0xsd592YB+CkU
YU0ACzk9aZAnbAacXxT2urQjeuzEZrtdpwRbBiGGs59JJvmjSMjY58omnCceeZVc3kJLy6akyWAr
kCTLUWRbvVXmiAkGu/+4WR10+l365pamfc6a4do9w3CPMoPvEQtuoZp5ZdO/aPiAGNSvEul5o7UM
BtNSnQAI6R4MFIaQ8ZreqJs+UFytKHBytWgJ2P4sVOmIWGTBwa4BxdU9CmD73VbsJL3aHvfvms1Y
J4oWknCpUjbCQ3WJ3hYc6kHKLKuc2hlsgv7WnZeIKZYeRoYklmQreng68aqICk4KKbiz8GTVEFOE
nLupWm2mGZdHG8j5SelS2vfc6PFMHlEoH5uMOwVGoXvptJWrZcaEaU4btk1M2LCKeAgNMqtNvs0b
lrl6MLglURZpE+WoRtIwphZUZzsSQqcvt+ggyeuvFmVqSqJU+xCBDKyPdHW/TR4IWdKvxLwm+0xe
ORICiF+ym7IoToCkUfMMYHMfpiQvDMVtGt0Vk1TeL++4Ow9hBfuuhZvlE0tCDYsiH/X+8GFZEpOT
eoncd5QZ/en74M8UgOvZX3UPkUfmAJNe6/Poo10NtrmWWvJ0oEaOKJDxoN9n0VqF7emQvokLjRl2
GAyy8phi7lO78Y38XoSxUmvSaWbrtZCfy+yBmz1emA50PAb2H/5zX5b1zqE0lvooKh8URxUPmSST
8vCXRMlqYoWREtgfRQWYrufdpvqphQR6/EK6zVdLIV+NPAiR9zHc/+mkOPEEl/rw/84orNIOZPqx
HBU4EG6wqQg6us6ck6l5h3LpiQDurcnEUbNTTAGwm9vQLa+ZuAzao8isPEvHPLJu98nTp87tlHCz
pvKNVX+GTAwbnkKnEdoSGGQkJKGKcG7aZk9TEiTc+C0CtI1XH1GvusLaRfDzMEEUC1Q/BvQgWz5P
S0RezxQgH/jYTK9Slu53d9ifmX/owFYF/MqL77dqakLpu2T+1RMLqV6cXV4bd2c6hEeXrOszSVgO
knHKxfClWWErnvU+aDfObcWjNMGYTEM7xjRRXhj7MjIhF31C2qH7G4HsacMI7mz55pgffui0/rQ/
02kpNIcY7tdBaO1LXKsIXD3wjYEcZAfB/LBxZPtS93dzElhwX7L8tlSyZU6epVUGOhyEqyB1F7G9
5fB6iQJ/6owRrF/rE66IkbhCYWL1QdHUbim2VS6/MOxh1n3+oxO0fPaEAtZpYTbVo1+QoH/+dU6Q
i97cuIuM7LkOWvWEjExCKWVqgRUj9uzutfeM0nw2CtytKKn5t+RLnxy53oEkxKF/MELlVqOBnJir
+AaWCu/TODxQ1bLzORjD+w5polAt+8umoGVGLfetKlscqmVwcWV4C+I60lcaueMFUnnuxrlBlZkE
kbAnnL23KfsR0wd0cdb/nApahm5k5SlGOJdTIMu3fcfZy8gkFKZG7NL2jayr3r7mt+8uklJaMs3M
AZtZ4VngzI/5DkdoaypIOcuZdzocuvL8HdGDNWDftiCdyCDRwf775NM7XdxZxYDJ029BtChGV6yu
1GDHPTJEeIW3DgMxxwra8WtJjL5+Yn3PVtMecJtqWd+fRhgSnA7ZKThwGdchW5caKTTxAFIAqzZz
2zL5Pea4tmMFfV1AdaPOX+uzPsgowoLio4VmRDmip3Z75my0fdOGLmezzfIyqwzR/1YkHWd6zMPT
XsFwJ4C7dF7ZHkTsrFPiiOl7hwDrpzaBccO2wPMK0QtHQjniYpQoESQ/J+wbgwIR0yeVuqU6rymy
NZvIy4qVea7ib62cpujVLElCqBjw8g6mwAWPlfpc0usRVc3XHq9EGhl0QpD17sodrD8rxVRlplhz
yp7rL0e2TQieBWqzJXbsgeuowV9a3LqL0gYE76H/vtEY5EnCOgDp7zqV7FZX4rZ59DCaKNFpkimG
1gFE2Qg4NPKJ+388pdq82717g388l3q1dgcLNczgR2ljSmBvjv81SWiQA1SSZ7307zFzvedMlMC+
1hwYQ2vPYtDiGZHZgMq+UcxZHcFvyopwT1jufZRgYbJBVJtjmEKnrpOrcXQSeP4PJDUlBgevKJ85
qJpD5YkaKtWqMmzztzSf1qEvl1cqsG5K/tuEj7Uji1sIcFv5Jx6JbnOdAVpWHrrE+3yDqwER79pK
1nFalumHUjArNly34mRAVXtgP1PwRfSK97JUhzrGDFv2aCT837o2miLzy2S0YXIac9hhpBNkwPlK
KALVrNDPvx7PG8esclacNyywj4ba7ALIWXIOd2CSdd79jdVhPXhLCESt/Zcyn4It/1HSi+NGitLg
SvFRDULQdTKmf7a7FHpmNjuwshPB9n/Yt9RY413gTGusl9SgPBySlPldKlQuw7u6BhSe25sQLE9Z
TkfaYhmeaISFgrYShuzgbwDt4hn2EaboWxYVgD1EAmC92+8Lv/UZ1oMJJPUiAEn26se5eWoFHaOe
XnIM2IQNkRJhrU5d6KQT0+g0E+qISmQsQFu+ZAMu1oy1/vKJaMs7cqDrBO4CJg8flkKHFgxXcXWH
kkT1dqzksyrG//owWUYvuLXlTMc/a+zn01coeb6Z3V8iPpz9jHE3d2N5d26ZEd8/VV0zQqLOJ5cw
QOs+BzVtKBjRNhf2HIq+/CNYWBCqjRfPf3m2uaKI2qw359o6SQnSl/GaeDRYqCiy2uOBIfs7+zR5
inT8jV3FfePRR7cZV9o3X8OQk5C3InqbwDJhgguMYZjq1eXSO96viWrXZo5ZoocUy8XaniL2PUVc
F8Pg+Te7JpmdNWWwHD0mXqBpkzPcKmN9xHWI3Xs9aPyyNrqjwfzpP5elHsWRAuvoM788nkLOO3LQ
eUumKRrw/sxJmfWgCvjGDDPlmKaZK0c1qnjJHl/TalK0dqA3+MR0CfgqUxuRsoGJSO1N2nEFSJuX
TbEuK4tIHj5eEfxnH9ItYlRQw1/VszOaouXkM86pNwvyUNGHCEWaEvnExTnDFWSFaKFowZ4vCOxk
bRfCEmu/02A3KllGiLPwHRdTBqjl1UyZIcUscKh/29uoFFebCbQT+JUohKTh8sI8a0NebRoHpQcL
1x+ZSEDZOz2FMUnDMYoO4dBW2enG6V+VTsxBldr2ms1Eriu6vW9+LGwIETNyfIsOGWRnKHmH9Cpc
dkQvyZ6oZSYtw9Fbl36bLWAXqq11ZAkUe3its+NCP875GlDSMdumq2f4wvynUcbhQEd9rgQxzL+c
COo244IQWC6enqIgPGU5M3ZnFgev77gzcTlYhysrwV29HNY2yNZCuypIpKzerpJl7OR6HdgSvXTc
HYi6CoVuObhUF1gNxzdLtnvHMfoSVs6I7Mgc27pBYy0vrRCEEGSgfdqmKKdSIw0Ohs4LudEHRxL1
tZh5d/mTlN9W036U6vqD+FN4fPmOIoFg43swby003oQx06V0/iHnYY+rOUzfbPOKJiKnUwtfxrWu
j9fic5lfaoOu3iN9T5mntiOZcgzEtuNHXi4ouxO8U7w+KezwQVrS31fSJgaJ1X0P6WGth0iiPiIu
3MVb6oLer7AblKn7uhipPAIsXvVNbrt6rYpfPCYZPnPBoteko8ZNAfdFWnuwjBYkNFf5SpXYZQog
yaWNS6P5OGQXPqzugzHfWf/rn2GSloWWr125oQjUknAX0V3p9IH4+JT8b7HzyJHsw+qpH1b2iycI
M2piHwHXYPdUGoSfyRu7gc3P5sxRqXMlquDxF/9HJruYJdyp3mkFXGZJSixNbDaxvTUWTKNnITQY
9Kc6pgvaR/3CDavT7k3A/2aWHa4yhj8Yf86tsSqlYUVkh4v2YWK5rV2D2eO7vOrYQBYsooywwMRw
sjvytrEtcrpYcHeRTdUNElsWAH/pDtIwuaVS+ZJQ+LL7ZHduaAFcvWqM71TjmsT8M7uPPutyvNFT
xVs2OyCOQWSoWzaNq3SVddMaHYnp8uT6O06Prqi8C1MRjODCgFk1TNwM0zsyuX3faWVWWcUqn8rc
zp2h1DozOFTbGuGcdYHUwOUDmp1leOVX+ngs3txm/MTUQPGXfeSlN7RWtHjHXOXNPo6Qz7S85D2R
BDMUrpZ/9NQTcYEtA+PsZmBl7Kc98crJXMlDJ7x6wVw8DBS4mGk6kvVH01bUeFyncuALXJ+eL8/t
saEzATi/QAy9tJFhT/jHGuw8cPGu2ltVjtAQEOcwN74h+tX3O1YvdKoby5ZMwwA5qmFidsY62Bqc
M33H8Ui1tpe8t/oUP52LCXOpuIgnPNLpgjDIBX4RDCddMzLGRhGRzLmAIcmWYAdPtJWgvX3kvki0
WY52Os8MNpO+upYBDWbXPxSOO1QHpbxvdn96BfZvWywf17rxpPmRiTDgv4TELKMoBlJaq6vNmjBa
+BNDd0ylSGOfvVaNXXyJt8r33Oh5XNzIGkhF9c+7NgDu87ndgcpNJTfUbabk7DqcxBmjtSBjzWew
hZXdY2Xvwib2yZSxNdwdstcQoyiAuj9Ieb8KyO8TMn16Pm4iX8Jjv8iC4L+fb0BEmhzyE/WctU5j
ZqPJa+Pu4n8jROBtmwJ4177ZDZVwu/ACpJymd32BkNpFVf5YlmmoI3WMUmBlDb25q9KPLNsmm1YO
0FsGVFlIMnqIfJJWyAiMZPHqDH5zS/KYZIFVH+hQUctWzMqHKLZgTVkQvdGLqlAa3N7bO3SAIAUA
cq96q/59zmtKYnp7udqnKRPsMTTJLvep0cgtAcoGCOaJmPxWq+49lRCH0o7lMQkb5DG2bZOT6dg6
Jj5v9ktrcz8AWtcuWmJNdjECgiEIyHqhdnr9HzQWD6YzZzdFCNxe1gOLtNXlNUP9b1MBNhjOwEwL
wooQQs7MSIjqgppauk2kqIWTUJeOcPo44yCTdGrKCMD3L1l5b7shMlxqA+KCQ/5ZXtoQHvldWxXW
clS14B21kiWcKDlv+cvDWnG4Q9gEXIhqAh6c4a66BQgpHRLlzgrexP3HaleBe7pKCe+s4BG4/zDZ
lbXAHVngGojKhB6d9k74Q5c1HbdaKxaMT4RfT7qYTpAWtepSTv72l/BXMVP/GeaIbCiPE2GXm0tY
/BmyQfbTjKMDEwmqOWv5FYsdn8K69vXVg4XtOmjpKJCfBm8ADKJigpa8NTVUvBD3tc4if7wiAp8s
9Qga5gyKF8HXZIYMiedG/d/A9+NkYPUm58vSlKdV3eckj/wfcv21VRSrBt4dxcf34ssCxaibId0/
G8CCGMCjyQzDyZoLIUAVpaLt6K7r32M7lJLioczEJwhBKDP2h2pwUun+69okA1FRKLiAU17HQ4UV
6bEyBTQks9sZiaxE+T3BGmFmJVqdy0qz7wOR7givxUkVlpaazuhevUDkuWLSWqEubMCYD28CHt6U
cT9hKnURyUAoO5zcTgLO0wAG18KQuSoX+FDUaf1mHIOUwq3kXeSrBpc/DsTKKE8p5GjbMxPU/6Mn
HdkzIPQYOWBkStRiW5tZ4/abxkYru5moxyX5sBzTKI0cqQQTf31cD+T5AlKyAVzMN53yRw5WQHNj
WYzpvvWffZBh4ihXiRiY57MOVoOX+FNgZ3ywu4/7NexmEkCz//5scEFc9Yqz+Q0LwzFKIFSXqtnN
xFzSgrnFLnLCZ7iwj6GIGMFevolY1Lvp1faVe9WEZp46xvgXjWGxMJxkLToT00oRIEHHbDQSB1zE
dQIyXbAcS4GEU0b3PIVckYv3aDAofxsG89cuM2zK8tYl6uQakhrZbu6At3jnOeWo3P9MXbTip+vO
WmkbfSu9ZpohP7R+SW8+mjdzU9yTsRsYLGpc3q1RfCJ7e2nXGNQDh7MhgZAJIigUcAt7yrOyt5hO
ZMd8mx/l4R466fSBn9/tCtqoa8ZKJMSRqXSRr8zYBgWurTZukkU6GKGf1WOafMpkRCUMXYC0I639
rXLehejemx4uNR9T94fO7iNRJBCHzfX+/tYishTlhv0DbPjJadKuQOmrE7YZLWP7U2b5tWaO57wI
AIX5izRbfPm/JSZvdjCFhhKVGGm5wsejQQ06v4/ykN4QC1DeoSpHDKYizKQxbDKOI4R+m1UFCCHO
EOJlFluv4j2y8gsswdWqqvWLxnZYyRbO2zUggTiF3IuBl37AIuiEbzR2DD8o1o2rPDJ9YSNS6xfC
Bz7xG0vEmtd4GPhP0WYBDci6jpVv30lRyM9HVf+YUIGB1vRfaTDEUQqLQhB76ZjqpTKvMxIowJGe
7XOhLiS9BgGelA3mYs4tCbTGYZJz9UznRgQ4YKp4UAoS8GKeKKHpr9yVe+Ff005nWerpGgzrgB14
mlnKjeDq2BE+EpFPwtVg87PvXwDHo43L4TJxkSnsYkOkS2WIJRC89jLN+JzbTfTwPdguqqlGndU4
2zdxrF/letbZLJszyRUrv1eYJQgk9MLhKwjz1YXTQlaBbXzeuT5gHcF9ubuQyhndfBDSKucZsAYX
Etr+nh+bGp2W5OQjQ1M2XdsO1xtWJtFkHs6pQBqYsYnIBtBz4faNyKba3+uis0VYB0tQbwvkCgfj
V1LHD/JygHMO3AnmaxG1Zt05RWZ7yU7b/rMl0JbgsgYx2bH7dW02oJ9WNWbpVKd5pdjp01tUPefQ
0x9qfDJSmxmTCBVrWURT+BD1fJbkjUYRyx+Xh6irm/lIbA1iDm3rP3eRojw5EekLoOTajtgTvxqV
SIOHhyhuffg+g3W2sfLuemmcYgWMXyne0hnY76aDAV0lQI4G4BMv3PpDC67hW8jcGtIBlM5khXDn
sN89XE9jlED/jo3d+UCsSOvwCk6a54X7ddytzl1Rs+gPpBwdHS1ab9zJkU4ogLq5YML9HZz7X3IB
/Gv901Hxoln2/NvTyLi/evSIFl8r7rDhIME1LQoLMJx+fu0+ZQiWjbb+pF6p1TKdCm2PYuyfKqTp
7Y9ErX8ioTaETFx+AhGclvKSkpebqnzrY1HX/n50zut49aW0jM+KiqQwHabrXNg5nCvzp1M89lPb
NZKOZxuzprO6s2Ljl3wSE/6aiL2mWmwd3tj3MNb5R2TpI6mdJBynrQzintCQ3Wk/t+68IuvTcDLj
SWE28CO5RcIZuJIEK1ypYWXCIfFBIAeFESTP9WAu9cGmiG2coiG8/Q2dL/pFtPr5bisWToaNCu+B
hfKKBi4YPjQUuaDsYjUmO8VGkCoPLwkwJWEjVtA9Uf0CJPq/52KkKMxnDgulw2o8ICWe3HPE6C4p
1HTn6J6V1Oq4b5hSvdzINbgcUsbH/msE13rF7Y3B+KX2RnnGZZc+AOaiGxE9MeNygYVo18wqPi0V
ZxVJn2bVXWDzGlGo7+ZnjgZ+ivF/XKgq5Cbv7P5MGJKcKNaNyeEZszrkVqHjiHYiXWaNpbF2FPPs
HwQInqtn1KtMM/5U8kLdFcvjMYvxx9/GY5o6XQvhDVw+ag2G6cKL2a90n2IWBzrv9eMpdoQcmVBF
LlGyy2ywKQRoEq0qcEiAmI+dxomRH4o/8/MQPgi4qpe43WlD9OuQH1zZMOVYwRImfsmQAXxN8xD5
8YesGjFFImuiIDYcZ9atiwCaoamNcfi98F2ISbJPvpgzoN/mASGE6BRcH7aqsJpIrQouKEccVMA8
FO9uRAvYn6W+cWjDe94kwoFbYOaa0NxTcidPrL+PF8qRSt0znU6Kf61SGqvTtIua6pVAiw8uVVRE
NMrAFz1vWB7V4ugAhytm1JcONTv7bAFr0WYR9chGoGe2ymyOH4HRcmrrfvXUqQ8RivoXZaRCsqan
Z9RH3EtCm6bhRqkzV09UOG/YaJmiRuMMGJtN8ZyxFUl6Y+Cy+0/UTTjfFLNjctqswX0JCFFkxRGV
HRR7NAIewlsAD2fReEBX13KVhHZIMv6AWspvlna05SIoAjp7kmAN97Sj6PT1rcUuwvS3fQU1fFJJ
Z2Bie+rmzkA7aKBCZcY42env3eOpBFRS4VeRLQISH5zU4on+Cqm+VhIOE+I/qgo3mslZXy2fqG8O
n4Iip51Kv6lhGdCAPuJvRdeYSOSkjxiVjJcTotccGhfyPgUlVh7f/nQaH1s4IafGG+rQ4VLPXABF
HrMDQi4S3aB7vP0Im7tCOc3uGm+TnACl1JkB/QdYniwuX37oaJVCN5/vAYUx1R7mM6zg1oEE+py1
2H4uH8LpB/iusgHbBgLwBB2UtIY6CuWXYIkb9/MobFpIvFuNbvtQiQ71PaJ/IyRk3qqv/W5IwoNJ
HJY/mjw1MvqG8I1CAICztCdhHWAZMD7r9p8akTc4dnjiJfuip+ep86S+3N2ae+Y2W2RTjNiNyX6s
3nzp0uEcr/4FjPLV0c9XSrbOQako8Wm8JKCKx+CRjYhEG8ENyxOsJfRpamg822WInsqXlHUV2E/X
aJexesP8ZGFyJNojnRMSld6ojaFYAfcrK1KTx16f9Yt7X8mEjWdWJxbjr6TExMDEU2wmqojcCn2A
lVDjjX22gm6A95th18f5sz2pvawEr9UCUZZwtVpGmKxJfSl7ORhuq1Ab9Htlbgz78MiYuQpbC+ed
Z5FCQSWRaCKucju97foMMmLRoxjo8xHhnf4LiEgKnSoq+IGORCAHs2jQDZMAWyWM1nRQLvk+YHHQ
TKGS/wXhvmBaDhds90ypkcqVGCrdsS+sxV4+zjnauNL3TK0ePjj8QcsNXBkgu7A5xgwGCl84kp3K
b255BXkoe0aVdZVf1oqJ9ufipCHUvyqv78b9FhUXT8fn5Qu0sOhAFFTnF2AVo2cZJZ1pqJNTl/nm
aDd4c/ts1/EpUQ07sv0NlbVndKJ0c6e/cW2ZL7UEku8xyzE1UkwK4+BV6BO4DgNYCTnyHKWYwyHR
KHv7InsRjAkA99ER8nprAFCfBhgT61dSz2JasmfyTlcJolf77T4jq+m4TzR/FBRc7Svx+wNHWHxp
BN0jmhtZDpSodn64vGAwpBFI8hiQkKKU3qvA8H5JVFLYCRX2tgrmi3K6CQFAgQOL/nzfJAQr3Zpi
QxLW+mC5yA+16HyvzqjkOAz0erRSK83R/gbvZk7Nhje7rXFBihKJitq0Z+98K9bUiNc1LVEEJPmd
v8YnEw3/7tShpS2pIMo5CawYWtnc/sgLpBG4wofsINDWZGrlZSWwzWPKxb4zr5mVRoKttorylsQm
2gOioc45k2Orglg/90YSJulL994iQ5ZvFEQsWXYoP+e+0NaT3TqXz0pZ7LCELrzARxKBqtMRTf8S
UenIr6S2vcf/zoCG2ylf2cZOteilFJwsYlaMmE2LjfB1uh2hWkTTGJUY7OxFjlYhNuzSji85CJpa
Qc1XUNOqOAF08A2qH79CMUgzSUYerPlgzFTHtmw4rmLrCd42LXnSwyto7Hq1OwImuiVytKstvTDR
deAPZE7kttM8m3y4zJJh2HN4JXlYatcLvM3D86xyRWaJ9oVs1hu37VnpWjlx/WaMIiMQk8ZaRFlT
VJhMBU4htm+EvUSb45X/beahJe685yG1Z/F/wNS8o4oIMsz5kkvEDeD6RjUoFpW0LW9XmeBtHHjv
J6rI0o9JZbEIqn1SQucUAJzXs3tHJtV9hYsQpAt0KBJT4JpVcyBQ32gh0KF10ciik/wyXGnguKZp
ZZPdzfgl0Hm0VRnbP+3ZgLUne2JkhgLJmuQ+/CxREjMqTU3s1mvDukco6Brj/PMcr950RBvSr9nx
JSOb5RwQStGKPyDVVO0I8Z5cXO4RgnMvWN20oS1+lPXUH8aTPf8TcHtonaYgKkX85udPCL7vmFbn
i5J8dwrmlWrPBzXwvH+CswOXMMwKkqL5S4JaT7OqIvRsH85BJ9fr8W5GYLr5mz53zzai4qx2/YXz
abrEYabtfVk+M9KRtR2QpAhxuHzmWGel+gY3RA4FBJvZ0op2+T4WeCpydgTG4qQIqPgW2LYUGYbt
pSwizlDScXGqgTxSeFnO30JlFaGrg7v1SBuNtFJ7vxjmmLHCUTk9coyiwGyffO8XnCP6SWOt5lNk
x/zW5Yz1vzyZS9TcEnUWe3Ap1m7serPETSAzdTm/YA/SihELnSbFHvTpqgzjEAxdOvoDNtWWq/9y
LUMOsmuxnVmsLReQhGgB4Igy0EGiUFp1WBNAk30jmcQNbj1QMk9oDk+JYSK87MNGgkUBT22SjIWM
Q7zga9FLIgGWDKgdvPgYxxqtw3IoU3LS6UhvnDaglbC7MczvmHDm2nyCcCABr6gCd62e7bgQkFqn
bWoLXmW9ou6OwyN5fRUTH6kwzAshBdKYcYmFYTUssihrGPrj0P2xC55WxajCWYQVh+EZ/YTrRq0t
MIzfCUr3KVxerZcN9P8vbfS1Kw32ydP2FI/jUv1RWnl/sCKgS1UH9/Mxm1RGMdk+9cB+vItR4R5j
epL7Ug/IEUe9ryPsMLNtuodvWqr7KQbQtyHdNz6gCCeDVR7iVtdiVEgJq2BqGQlIqfSL8ZLjxyM1
7a8xH23Dus4HPJw+JHZGSXmaQL39TtGLb1VP6smUUaXH27CqoSXF7O0ajUElbqWR+h6Ad32ZHGEq
5etJZK3rw0ImnEHvOUAb5i3BIN5oPhdSyU+CI7fhgE8DM9tipENUCuTSVhLJFbFXsqkglfVF9vrF
atmA4hsddSp8k+E8AVz+pcK4ZO3NnHIiVqj4y5LnF6qhwf4AXuIdAZj8VNxjJAoxApVGME92UH5u
kir3IDe8ydR8/eZiP+mZUBwdOQdM3f1DI7UrGbTuAkeAotU0OBKcDb6VSWIyR6UCai2dU6kzU/eu
xCkHl5/GfzdzyVJ440fTqS/2nlAVavrTv0IDW8WtH/+BbcdiOiFhj3hZAumhzG/kiTgg2MIPUeQn
xzpdVJbzgrobbR2XvK/5SoQKfb+bBrnrFmgMO+KWmDlL262wwEj2h0z1vcz40IL9iFzAfEP3hReO
dX/fHSw8hGFr2OvefqRTQbRldEhFSg6wqN8jZTv7j7mqu98s3zBXcguXV0tsK0SwVCTiXuksDGKj
RiBAki/EptVnorvYoxOzK0yttJt+nNucsbFXjH7oO+4Av7GKbbhBBcE6QyUnx3vgNj1NDwUGHlGF
r44CuUj3C1hgdZsDuC63Gh84q/bGqN6ZLDn45Bn6x+iwxCp8wO8naLW53q5TTMU5aS63eH6b95jg
eHIEE8yaNW9+kgAE5p14/4eNTX4yYI5TtjIHZwNMtuJNUVV4lUp1Z7aWv0Ge3TR3qoYVXs0Gh+Gm
tPwrH2nT7c9V+QQqgBNuHwGINqMC748UfHAutiUXUIDgTo9Z+GsaoBtFkrkLfdB8ZqUik17PMe9P
LyoDzZ0l3Aoq/tzHYAOdtswy/ly81ULBIZrdr8s5s8vqaN4mUMmykLX/wfZFVXx757CK9665tOzg
qwQdrz5Y6akcHJbw+d3lmCRby2Fzoi3Rpzq2+4pFK/4zv+8hqlUqQ0nKGajZSQTee8pFO4DLwjXN
Pd4/2CXjwufi0M0LPfED4w5Zy4Evo59nfbLqBIw3HwG+YhJLE7z2u9Sbq5RlQnjynR/7UllTgPfF
FrBfshN/1ivQbQoZ7ODsoHH2znmpFb06aAqB5Mhg2nrsWVRx8hOohMLxSlfFlTwgK5DZDXJ+49lx
bimk/dtgvwJaaqWly68VB5JVFRTBn6Wi2gc5ASSEE63A+6C6Y1b12F3GRIu60x/gK64HpaeFPwY/
9Rw3DwvvIWtLtpOylvv+CrM+/kG0lORmTx7q+PtmbVqbfyB0MAgGgy0bs7Yog3+DA4jAaFf5eYKY
zphTfiMVsUA3/jxkGxdFZ2WABgG9tMdx5fu4xbR0VylnfkIjefHz7i7opXoDvjQoPSOhQ0z4WMWf
jUZkh+PYf4PKcPcqEeJnCON7yfCica+XmxQ/Ksaw9E2Qvz0HprqCYTyEr+j18jaE3gDwAm4G1IAl
mPUD0n4l8zz6VvmYcwIk0qHLrWG/LFiFGdjgQcsxQerUc3iJkOgHjPhegcXB3xA9VgqJOj6EOMtL
9YJQFDaaMfwXg5Ws4pAcaUaAi6iMr6Vwf2EbslxQ/UXFDq1Fp1QmQK/tjcdetEcGkD/tRDqzezQ8
MkWQSBa9goKaEdCY1YMVS8PTc4OxjxOXIMg025opBtlKmI9Emss/Xkbbzu+PXpSzSyuGk+VCdDOp
VwgqbyF639xVd6IP9iaNOXLJwAUXvH0r1RqgWsPt1eMYHQAPysH/FF1uA5qaKzYiIRByWfwK0kfp
ZWUS3eNZ4+zqa7CYbod4SaxPKhknifRy99TRBDqS+CdFxvzLarZ256HtFVcam4993H66fTpeh3qs
39RnzNLpgPN2SrtRQ3N82Wa22b3xsNRYWelwH69dv7T8H56N90911s9xQZm9mIao0bqoGdPf/6zV
T0GeZ6HS4Sp9pIYHWT8+vIVlwYExPEewEz2xaYCmqT4GA9KVDdKXK9CXw1ZfDgS1LVKUpTOnn1as
WHMeYBkoI8py4LdUSUgFcfhlb3DeSPCNXvTr155yE0zyEtumwhte+fD8mJN+tlIT5GSw/ycxe0wS
882T+JNocXOTqtiRVrJy3sCqiEX42fB6eA4K7d63K90VN7UPWfOYQKLG5lWH17dG4A40bdgkenrD
zwa/Zh42NvUNfu+Vi6zZ5QG9UKKwz06WzTGvms6kHh5KM3oCdMegyrQN0rxA5pet7vJPdWOlq7gH
TYfU/d1yXEH3L70otygBQh/cE912mYFa69fMmR7iTpuAGeOShBPfSjEwRwO03+fAs9QfXjJ6cnB4
bEHi3+5Yl2R9mGrVA33wqQsJnBxjGTucOGYFYhZ8odjT8yVevkU3jdk3GcRjmTSxzHjXvoOGTELp
dZIVHlKHt+Ld+RhKBCx3mMwT3F5GNAYiYJ7UB5QFPrQc8Qde+nO4Jap3PPrQOuKND8AY4ztctYD5
BDgo/wErzooG0odPXnlE26n9KirXOxUzzNvNk9WJXUGqCAF05P11nf6FzbT9IiSin+BSS8GQEjah
x0xz3kF3WO07Z5YeVHYVZoP2k3AA5TUCZRiDtA662T/U62seJ9WT4JN+0JwgdLArc1nFDNyLQqqU
lYknA/w/87WaQPz1DU0o478lLbDfeDv+nf5dVmihb5uaxfpwrU9olKqhLyI61l4WN8kXBAiZPJoO
icsJEiLNoSgMzfSoFawRMd5oCBJEDfxRbXSFwWXdc+YFp/iuOFuo9fr7soAiq1XzZXBjaOUHhxSy
xQnKQr9zvytZNgd1x4u15Bi8Q0zVExMmScpW/EO/4+TjuM+lLz/e6ALKy0YhrH1uhD6eM7sj6SNE
IW3Ta5Ib0nnRcy5VH4x9KK9NuJGAuBo41Xb3o/vHb5VHzytiLv7Ii+1tOFot8dMR6At8/UvtZeVB
fwj8HdFR8FLZ2yeNCmaxNTEnC7iwhjGUL9pOK2Q3787U/4VwWnC5gnG3MnIrslGsn+Y+Kghj5vvr
jLH4Pd5b9OfdQ7mqYCaWQOnfwxUXDPpOUK17pCq1s5JiOLDmpgtTY/2a3V/2SsxqzX2Zo2LAqHZ8
U67Nd8oIZ/xXnmH2yOTIkQelp8FyI3PwNvdcvA952M6HgdPxl5ctD0prLYrOGVceSOHK7xHOQFAT
rY01/dPxM+NcF5PoNjJie5gvwsiV9/gvGwgXCmf9hG/pEiYUOZV2pmUVwvSEePUydDl9mc+I84hq
P82NRKMMcvEVkHDzKJ0z/bkk3QJQ9hWHwGPVfxx1dIKvRN2laObn98NeemrJhqgm5KETXE9kjdZL
FCcbu/2d1+G/cd3kM2pY+5JhdAJ+8T7bHmoCfF7F2KF0FDBd6GsAvr04LKluN7PUhFHDoW3tRh1F
BJWP+n7M8dUMf2Ueijcc+FkmvsJqxVVg7QlB1N8lPa71QNzPNlg1DkYdRA08Y9iTikLbHoH8J9nE
EcN1mApGSf1Kxy97uicYIlzUmJvB0AsHsrxoROEzrNcKf2hoKUx0+m3P5/HqN6TmskTNvLwzKYFn
JV3ilIISOeP1LhqmppJFqPpRzAjs3nrIuLmfbATbprXdgZGbuiU58L/5wSaQIxkC8oWR6PFHz5DK
7iw0Xv1/7NOJpToHbMC4+MjXlUXc8e5GyyPNH/cR+YYAve/x08y9baGOl6fdDwLc9vByrOfgYQ1P
z3xzppX5ZZdIE4e+x0Hs67MGveYbP6CzlCnpk9fcgxAIeno6gAcaoNXnRf0K5KZi0yXn801pRd/I
oQaiGx6h5BC6LOmc6GF1bY08uc9+QWJ4U+K4byxZ8CDrY58jsciDSaKBVge0OjD3i0hHRtCShBg9
4ahNGhKMl/negQpX2wlfbMZGZzcYPBePmwuAbWx7fq06P9vr0pLiBLoYqwnoT76B2fqnNbk10FKW
dHNoHJ97PX8IMiE+3K2/R1P7p0k51Sjfzlo0UBvdpOs5eWeRme8+lPJ6xjW0nCnNfJgV5CrkBc7p
qiY1mgNm6jpNJ59jldfDzk/rluYRLY4ANuooFoNd7EXH8u43NfUaOrhVqm4V3/halUOgPB9Wrkrk
m6SuYcpgJHd+QNG5Y8PeRn7eCJMis+yWxNsDzhrOjLL0hpVG/ncBL9YNsnAZsT/RXu5jvwjvLf7U
jh2T+DQkiJlBrU2t48gA8sFVerIh45OXNOZqTY/WYYRv9u2VZjicznbrNOf7LVMWiuhEAWpCoEcM
RZRMAhlmETlJiIGACG16KWAALPSB3+T4hbKA2fUV2GggXGyNsxyryrEhlYROAk8GS8WT+sN1Qv8t
Ik+uiKhMW/S+B9uRkv+6Sw2cT7cNMjBHhsWkRdfaINTcF+3h6jnAtzKQZit/7ziq87f4ya5gTwZf
b1bQR/DjP9zjluj+hE72AuidAXkUZlA/GN9701WEj0sFPJzjZp3RsfFz6QL27LH/dlVnFjD+RnCZ
WR6y0lLmmSXXDOF0PmAdVepfsK0BNRHxLUtXjP3SVrCT3pBw2ZrpM/KopiONr9K4+R8oGlGkYtiS
/o8K8P2eb7c4eZX2PdXXcVRzOgpSdMyZyBPNSl+yVUkhkArMU12wd4d2rRYDEQ12K7gXU9Pbofdw
zkZq/JDy8zJTbTASgbyRChK2FlfscqLO5z6aokmPRSoxabyBy32MobXrO8RJgX52Rboal6+HXDoO
eMJrE9JpIPWzvqa6SVxlCAbbO3zsFMJ9bZrvgDS2rFnXPJi59+TNSltE9N40omJKa2l7doKuxenx
2BwHOAP9EsyTTQgo12n4K31EOhWACCIHVvOeUd1FvZg+korDSC8qt1rKBBEYDWS6oDYWA/vB4Fw4
/UA7dyKKhEWXCGe2H07VOwWuQtSpY3AQp65e8x2vVk/j0iYwZJSLn8/uWTjZyKNG9Y+RbzAbngyX
RLaua/Rx8RVYrhJXHYyfiTuV9kLe1pZpukoVMg1FHX2P17U+IjCBPe11a+ow9+QEmZBCMVKc4rTm
jVIjYaBRU5MaeB/IJvKIex/mZja2w+0RehFqnU57LVKmL6lv6LQQWThR2+Am1yhMz423owymQ9/L
5NCnVYsgRQmCxdDgxqRmQAv2kwz3lzH+2DP4uPBAS8ZZT9mv8YKxgGNm6MZok/0SQi+iJ4mSIrcc
dRtf11VuG1+IzG3/cEBXXrxA2M2MvCIcDE+B2P0JCzgvkndk2IKq+1Om7Ms6FVpsagaRXmtwpM2n
x5pr5CggiYuv4XpTsnEzAK+FmV93wKVg2AoCDcRcW13oY+O57itbdluMODp+wNFiME1yZBeOVduH
2VfHADIoT9+fpJtjK/gpNnQ7++S4O1V3W2VxJNf8PBEJnBOkO0V6pipH+MXGk9ks4tC3/yr5trgN
VpbF3gAxKRyuiW6swStMiDfkoS/Oxr8xsotfvhALYu7AnCEOF3tTTW0bNYuJk8bIdjYZCD7B4JqZ
1Sjfkuq6CA+tIGr+9k0HT5bcLIKeEqUM0q3rAqlchmHP+zRYb/y+q+0TZ/bTOnKdqJXS+H4mKH+k
MuXrizuTWI38IMGSkJfzUe04Lg3eyBQwbf0ox+M+c8hlgwYGVIJZtNGgIEtsYZI5Iqalvei0d6co
g5Bilbc4p0sOrZO6kTyUTxR1ZAgM93xC2Lwn5FauhCFaMYkG7LXlimSJB/Ui77vGhpOEK3WfUZfG
c/pEX3WEgBcxGjKlh+YzMHmgah/D5nEYcZPa+JOkccYbpPicMZCy3y8ojfQepqXaKR0b9VHwlmsK
LSN4BzZPiuMgTvRTuVzxnGkctAWtY70z+eQ2chVoaUnzf8LSfzUr4MOWbOcZZ0Fd7H97btCUnDv0
bIYnUJZFPiaojmzlTlcpvZLvELyqbPtLxjz3hPMIK555EQh6elUGyUsIngiD1FXSjQ9vN18HpcHY
a2m1yk+WbRWWQSDjTdeqelrge3/gnrB3aZi99NmF9LjGiGz6KQJdaTxcBVbvLxosAOKD9xTVRFkq
x8qqItImXFRhX/nIlqULZHRjRBiNe6JsFISoo3E36wZrTRCYfRd1pY4kYXfWC8y47vz31fkK5q49
GUEo0VDc74709X5dn33c0QlvqVCA5Gdi6/GP1XJhJNyvB6KxlTDy2cgy7yH4yicdfJv0ysBFbMPD
oJmGNm8t71t1VocWD0zdBKjIP0pcTT+xlwxI6QZzw7R5aMydWgQYUVrF8sE2GUCcUxQNuYot6Py1
LNNLweXloq651Km7Hi3SbADCGbJyUpYkPwp06NvasRAp0p9IiNp4z5XG/NJMlcoXGmxwz2HhEiLy
jphZngJzCLyVe94tl23GXsqhiZ39tuNovrZ7/iYx+s+3m+EHTbHmMQyUn6AujHZpCHm1FMhaeTaV
gOn5aUHJ+GQxhbtOnEqhP7wfzlhzRacniuueP5PuKqeU5H9k05hoi537o9yLR82wpgZYnTVAYen2
7NEbu+ZtAxs27sU/IdZBz1E/CrZNdTA8aBG2wvO1rROUbogCfL8aSspuv+5VWCH2n0h1hIjSj2MF
ZUqRd3Wt5y8XR61UUROrvW3tjgRZbtDJVeDHqibpdE4RK5BF5hjc4yxd3TcEW1bnKlM/D/YAF+6L
ei6+dMlnLUjuSBt0h7gjjMf3FpcsRdhCfq2ny9kkMfWQWlw0bipuAIgMHdFZoyCRjVfk6fpQxc7C
hrV3S/8g8bNHkInFXkPUg90nX6gchXVtouzVtFhYmMLp0YypO3jd/mBacQiym5rWEGh4VIU/4fBA
aOVQjXklqk86KpPhUP+uS7tZpfXZpy9z7F8EMxnrKYAyhgpyFhJ1sZ1H5/Fv0Y89ipzSlriKAHNC
P1iFQcifMPaQHwmdScu6Ta92DjB7dGawAXxf/Mcgopksb/ohP1jE7j7eZWRwvW/LMP1oGNRiqYsB
W5JTzcxVsDWYuzZf7qRVfBMld0XOgmiil/d+XLsGN+HEySABXuT3psukbBbyFDwR+bd+WMaUyh3m
Y62MyrjCk5Ed95OlWt4qS4Uwuq076Fo6pDfN5/PMdfAJG4LNFsBynkQhwqIPOCKHftf7myZuijto
klJeEMxzAIgUgnI+uTRahnl9bhpYhzA2GTfEI1TqjmLUvaXjuF568QGrQyuqvmJCsaVs0ZXCiIuj
y8QzbMKfqP1KoUqIeuo081EE0BTqnaGmqI5uY9qSJ2Wdsb59ns78P++lUNunfY3vHdC5ZM9vFuuO
PUPi5yjx0L2UtIAAVvvLSxvvk851EQIIRLse9SOcsG0YuUO/CsbnPwb5YW0D3kPjjtFIoDtXF0i+
1Cc8HWY9tTejyHx5amENANj8Vijm3j+FqWP9AWVKmwusZXJllQkjfUn1xegZM6H0xEW+g4R/X6c5
Q2BH/qQv931XXPt9VKogR+Am/1MkAxlSbwH2pOjKHgqWEmmml20Da0gXIw3vIGs93z9Vjv6cZBia
crgJh8mzhGhU0STIWgHntc8L3A6NeFTc01g88SFVrDsgXISxdG8G7pgcevUIF5JCNalmw1YCxBH+
A6m9965GJwCPe3ZRD2nBlBMvpKwzcrAOM+fjvQp4LlBshJH77ZILWZWw2ZssIZ0MI6GiLUh0aSjr
WsGyzZK+QUwJo21CNd4soeqi8b+PlE/RAkIsUUUY73bWZHtVQ33+ocRy/qsw7x1I92yGBt8A9O65
nA7+e82QRv8xbUQ3e+6857y2j/fJVFdOEjjrB3blp8JtJ8MF7Fbu4lhNgctFMt8dflxJ7bNaVygE
4OiC1wtAPi2leKMFpqhqdX/XXP6fK/yDP+d23BrsG8XZfnIN3tYlRWN60Mp9169WQU/WNxucztgd
DsR0xePjfA9rmS/0g0rLunnMEDh4g5I3dZqBHv4cguRjeiH/NHebwm0V3uYGALotUFSoZoEVnaQo
mItmj4sZcS/2JPXq+G57aySY5jvXNz/uC7/pgzLkXyQ771qLsQkLiRoPveqHu5cpMZEjvUZc3axA
MlQaRJfujR2wE4bV0/ML1FFKQgdQaVHpCwwR9sr+iuFsTuhN2b1ZsWY5vJBZTTZ+p3FWq8pl41ZQ
eef+4S/Efi0uoRx9coMKqWaQw1wt++UEsrhKNtIDNCUzPVVnXGw6EE8510h1J+fy8rWzs0J93Co7
BHEW4SpJl7fHOELiw9ff6B+qY5Rbo1EHcWLnMqO+j+1GiG5G4GoDnHj+7Ld4E1WnkKVPb30bW7Tb
SnhrcxllKHDKWugSTALdah2ts6q1yKxA035kOpk2fazxADvEJnu4JxgwREhlGEtn95dg93ZkLYXU
R2oO6ShsO6AbJTEmEqiqLkmSyFjchrnG5mIZRHCIF4IgXlTTTjuM0DTVsA8/soukfTQoE+mSLOtf
eDh/ckFN+WB0HPdvfXd5jT58XafKfSAZfWrqVkwXNleLEt3CVaWf/1NfU4Z2CeI2jQS/7P+SJNQk
5Q8SnuI3rizc0pZQpFBZkvDVe67VrMb4ny7/QmhfIXsPYxubiozBAi1+9ugRNhnAQJFIJC0GQ76P
y71yg1RaklNho1PPiH35ApoPoMmkgapt2z9CQADcE69HAapaPd50em40WF3ynd/OHF/XuL7Nennx
Li2Jz6pZ7S7tzrNCj2+4XMMXpKegGe4kxZy5igzqnL+xHMEj1t2MEQEl8vYaKZE9+JvDCtai5si9
OejlE4kide3qPOOae7zAryHfkU64VJSeGK3P2bvxTccSqoG18WRKIDGM1cu3SyFqKzWoJt8PQmbz
cqfVYdz17iB+ndOdMgW8BQiSEqJ/Rda25qiw72nK6gdEJSvUIjhd0YX4m/hrG+ZMT3QVYukVqmnZ
fOyDS3TclRka/zUutzKbUcbaT0Dvq73MNpjdXxdFvsTrzSqd7+rS9ZPf7KhPNIj9Emvs/M2J4C7n
SpGQQSZHlMYB+Ar94yMvqJlsN7OM5sewFmUjZXNsxnC0oH26Z9xGc1hdcpY0OvAiZLAASFG8jj5p
rtRsp27Pw1OuqlB0lcaYjBuHRNka4as1I8O+T9I9yLlX8hauCKtsmm460O+svJgXjypem1nmbnuA
6EMHzr4ZA4rE8/oVuAgKv1wPlQoiK6EoFvwa8DpgQ+C+RgQESgb/6UGuLS3DJdWbfFzuPDvDkCDd
tA2NiYULmlGwOSuTzKSry9x8RjZ/PeShpkUkEmqFEgyApr6XLTc6LrBvGsx90wwYVVDC2C87489M
7VdTGO9Fy9NsKKdln6EHf1nOHU3GCZt0pi45rxRlZ+gghbTwCGGreD9spfry6zmXv7zvw6hSVRT4
upgzGvasxRzHF3j7N4Zh/xm3XRIYYpDzHe+4VouZa5E0umeUq6iv9SRSTbwG9f1Zp4oYdNOwvidx
b6boPE7ZCTstfNT2woUiDgxF1+xOHTyclervI+gxAc4oESZoAt8eZ6nki5mcRhZ/8D9X4WP91uTK
5womKins8NsrWpaaOJyprD4DlqXpYz132MICzUQfdAZpwXGmA+YJYQilr/Q0fTojU9/Qai0whM2w
GxsamMzKbNfdC4bgBGzyCCY6PCL4ujbPgYMA3tB1/vFJNnh4vIRpx6AmwykooHwsbW1ZUKgDJeHu
7O3vBv63roqkErWbYXfGgFHwriA5M6wBSULVxNcOLueP0czPauooc3+lD7QQnqY2VVt9PMj2xk2L
ODEECx802YkVxTgiOLDzPqk+shFH0e5teAT999JKFgDcpQNKjkuiJvGJPxhOUANvkyC2Dgszvjxo
mXtuOL7HiK/1dy3sKFjoGYHAfln4EZWVafIyG0xG+WhukFkP6Rd0dK/a+I+BawR7MTrArumyf6Xi
X7Lac6HJQ2K8JoPtCakuXaAOrPFzEJ3jUVO7QFRTbyMP8nE6heHUPdqTZBVDZwwjKhDoFaasSG6z
vxlecjcC767eInkcdbUKUkITGZPQftrQs+QuuBLNjUdz5rKZTm+NxJ8CMWtqbQnGtWTj5RPs6q08
MsKle7rsm4om0Iar9CUhJFzyEVwoMuMWZytNfRlWfIvYOkVtMDHa0ipW3WCwzhZ4xalT9Gf3oznR
lx7TieiPMB/eqECy0rRdrV0C5+ZRA+NNLIABPjH0CNrJjzTvGJ7Z3luNq0P/ouZ0A0Z+wXP0+RQt
Xq/q4iU2DE9jdMY9rP38mcpoIhqZ9M6HSWbz8R1+JHED0HrRrOunI6XFb8dg1+3g5+nM3qnX3fOr
scbMpkATengbphI+xGCqawIFtmElsseBuOVmSr95cg9uPMV53SceU6OEfu6o0Qs/EUnfVfF21s/E
KlJzK84Ug3JXnuAgJ6Wply4NisN6WN0ZMgFnO4vwOR2de1Vje55kQpu+9oB9sP6Xjc2pdGjDPDQb
cCXlea1tllIcwTKn/GnwNTklWhax+H8nlrXyalpAuIqt6SJ/llNWBXXY3WIQvIdIxBvajwvSGbJe
3mHYQjcI8ZHd0L7RwE3oCP/76YhmvBbPAxD/BP8CrQ0SvjI9yTTJjag6hR8fgZ3sLylwCYdfeaTq
gV9uNyst3/AZ2c7kOx/8CdDmkMwcn3j+boVGvbNUTsgubV1+xegxgtvwMhpkmELorSt/UpvWdAsu
srbiDUXMDQObtOwq+fasM8OCnq/MSWw82dFB1Jfrt6T3tTk9TJMnA+DpR0L0R42ExLCU1EHTl+sP
KfGFytH35I+wAXQuiFstl/OFBZgpa53L6r6zdzaMzguZXA98tdqESCq11/Gxg0VQRVvjaU/wGUQ8
h70HPtgMhO0rmtFzPZfMb8BrBENxoOxXuwrBNMSEW3iCbn4E/0zjGsdad05QeQ/y7nonrRCS4gG+
qLIREH2YjIH1NH9f6cwzfZxnNCTIVeIGRv/+b/lVnbn89lf4qUHDs151DEC8e7Q0xSzu2zt6OaaM
+17otlEgkvArAvy5egEwx44KJQ9h5KDpbm5u4II9OQbIH5batvCS4IV93Smdi9dkc3ONsflayglA
UYJNlpYoq+uplKVtS2LHStm4gGJukquCsiZJbjxFsvGAV2sehITEotaQKLSQ9x5fIQrggIJXjGEE
mfLHxBkReSPwUwXa8F0h1KHKSJ19bme/hICm96J7WAp3A6zuqwz2B5sIM9I+RFo5sYjvhdkbOpMw
VJPhBT7vrLltako4nem2y9kP/IWJJQI0g3ymzqXnzX2onvJedxvhOrqT+0/tl48oK0sBdCAI3x/n
sxb3jZ+qYZpM5IKGswsoo5AV8hwwxwC+7eNUi7jl0Gix/unKI9935T7JZP7gkClWat7WYBkFqd2y
Yg0SgvieMvpiM3VXK+LN6Bq7Olymn9YAh+QXqkTBKapsERDpqlrQ6Wk9SEOb1tfC5NViFQeu3uNV
orJS85LiJczYddMFrX/uFwdkiyiKqtwT6jOyFC1TMmbx0iy5r29uC/8DUpwzt4bXKvUBgUkbxGb4
CuO8UpTfDZkVMFPr3IERQ4zNUyIySDVpDwGvZodrhIhPY7vHk/eiF5MiwaqdkszlCM5UzhFsLiGR
jHJTvA2riwzhhZjBphmNL1QVKpak9IIuMof2wevetwosr1Lfp9egLlcAAlMJEcdKdAuluUnvFdIH
NpAjHfOde3Pa5lZzL4QvKFuExq8KaoDx1yKMyDZVCzCPqmKmzofaoLJGWakqjUp36BRmXYDBHPU/
ji8WNroTHAkash58XZZ2aTCedA/5Icbf/mmoTp0YpvrNn0xB3+lHdPKi+Txqq4aOFzPLqPNFUuB0
5DqXcI+UPTK0zTZxpR9YuVMa2BqLgVSN/Ae/U9wLs1TyAuaq0GSoUAY0xjn5rLNbaYsDJY/TpZ9A
6Y0MguZh9HXejYXwvLAMdZGDsyKyHLiyK3j0a0H3iN+Ojaj69v+2KkLLftdtPzEmrjzq+5oXfe9Q
zq8iKRAR/8Z5B//iTY1I8RLGJHDoTje3JvDYQFD3aNBMm5AfQampHEHfRScUakqv7jctL+kblHj5
IcfUwIL2YPcJwidOhcNONyi76FklNf6/89ystQr0s9s7UPxV4ayjpv26rPLwIdWAZQCAqZkuVpZT
o3uc84IsVGnLlOyN/DFaS/EfAALBBNVy0ZsOXx4S3Ta4T/BwaNlNKqxxDpwoOSnHBlpqBZOqS66y
OO3o+wWagFjhwEiACXRjJaUZwHseGtEgYYPK5CQFTuwca8Mo5YPNoDaBkQw6BfopZhcpcMJpyjBm
SXKgM+oAB32rM9yJxzmmJ+uauo0ppykHLfKw5qlVtcKKp9YQuqtdOyk37OfgM6PoZ3mcAISE1ama
W74z1nSV0KfJQuaJv1wXOkZv8aFolUZL9Vg264Q+6AhMzoErGESNlhbxLFcHitVarYPApFn99RGe
eDYopFp4y5aDzglM71Hn2D/UoY4bOvekojf8XwMYuMjQKRFIn2Im20mDwyGKy3K7/Jdwh2m/Jpc4
sZfV76PlwSVmw2o4hJgy7/d/okwkJyNuZQfLpUBfQWdomyX7eL4yY5wMvRZjk86TTRsIx/GJ2NEg
snnczLldAEUVPxuE6//Pp9fOM21vBEBvYoP2ZOyvpcHRFo0/+GuLE6534JYxD9XI9eTfHfPL3J3q
Qr5v4juEo7uc+3HFhye/zMIEgu9HVKAy4M58BhjEZ/V07BlrYv2M143fPhhcLXob5+MQomta2AVS
KZor+FEU2zKPyQe1gbeJ9mJxecIwwB8rBVFobRrNN5NwJg9/Ci125MZuK8fkmLSwBvy1pbWexFc5
JxBqVJBn2GkYNl+sJ8XurWwpnC2OSNEUJC6iKeZK/+Il84YSeHLvZ8fJSWhHxeVgsIgZ+7jN1t9k
bBjpDrT1AmViXmQP3haI3Vyaa21ZfXyYKWZo1GHDloVG0gNNJE65HYpKtU5BZylSFeDMLFlaltEF
md1r2OcHM4TEHyaCkWL6DYlDXRXGqbbZweTtmKx6RQlyRzJhqfzLQD4WP740UyN8FiPi2H3EP/8E
88CBBLp0hvez2WYUddpRWSPYd88cs62Y9D7HY2xwd4vdWRMxw1B7vs/EU5JJn3wDOHAQq1JIYhBB
nE4/ielLdC0FhLna8w4QGHiH3N6WwsztVsL3KhbtOSTckUbtXU+ALTbHoJFR6YjvUGgRJ/bnxhsu
n+UkXXkd8TlI1uR8ZISNRDAj29ogmtOB8uZ1p7073Sn9nj6mhrifuoUqxi7pLfYJrqSMcbd3ID2+
R3gue/jJpbeOs2XWVCd9N1/25rJ+aMIZhgGZ4M+NNcnmapK+6b4UWPH6BlMrcxYSsafusa40d72w
2ZOmNqUZV+z2eNuyArwOebuyUYuyj+WgslphzEHvHcFKvC7dwAUTG3uJFypMSqZUz8O9qAqUbPXT
megSQ3nFKXJB7xmxIysTRrWdAz8sUNw5tUHkJdACSv4aqxi6pp35rcV7y3UDYbTV+YqrXXMO8WMx
ODBCULmuyytpnKvPzJo4dYCAy3X64aKlPyoXzLtiauXK0lNkzxcA0kbPHjVWfqD4IlTdGzpOrIHr
93CEH9pMrMvLmw5P9tTms+83c6NCJJzxg5o21YjbehMaxT/2gTTO5XvLGhMaDzPlXd654Z+WZY0L
WjtWlbiBmNKL8F5W8dS+xZVloVarFf+lrG/aBk6fb9q9AkO9XxvCI7U51zmpVYKaZHw0ud185Pya
PIg6/A+Iza5J9fUcBq09Cvy/qMZT8QL5Dl9rIwyEJECL5eA9ANOXN7/7qLTCT5Ixh+Q4b5g7tl0p
9wf1luFEQC+wvp9Mw8cyouSYLmHf1LbncqYk2SzY/W3YhH5R3iyoYH90uxT//oXZVizAZ2WQnJQA
PYv7UPdH+aje7l0LYIn2h8QwZQnJoES0gGcxuxfue/4ZjoJdhIaP5yAmE4qV5+3YLTb+oIj7h8KC
BXdtVj4Ly5rWSJ5DsL2wu6Qs08eeCLqkfRxeF88PTBs8UZFceVWYjMx3hN17GggqJkRaqdTlQs2s
0DodEYHZVGT9xvG306cQxe5RVIya/dlKfwlmnb8YFHkqtMvk/AFxCNw8Mmxsdp3M7StZQcgjbVlF
hRsh+qPSeze7JLS5I4tNDUIOzk2WMg2Sh0PWC6v36WelV2DQZzxheKVZDxUiBcSpHFTxpZ0jMWtU
Yw5uzIzHlmZ6k9ItlFwtERqx2YlAdpJdTW5CBw1Mr6BzKAJCROE075z/WCcJS2h64y9W15EEbttc
iTDQ9nspprQlSNYV7+K6Bj1gf4x00TXTPH9UOY4pjuSMEZ2/gY2dsGMHmd4p3DRrAfz4j4ZP7Hx1
pNRm9RYCQX2I0z4hAJc6VWVCtOZ2xUZVZGPO8o3jN8oB2mAmaUdgMsqHqf1DbW6Kzfmv3UN1P+ay
WX7rq+YPlngAMC7wrghwtdJGUok6WUdvyHuLYBWUKi1Mf2aKiFafTh2Uvt4wXmZdg3M1gkyzonbj
MFPYSwXMNfl0c3DtMic0Xng47oy5s6cS52ncuDCS6JiZGdrm86WCzs4+7udmcqAqmKKKA9nTtNd5
zVY7tdx8sncoHWYAedieXqM9k7RJZVStopkgsOY3Twx9LrFsPkr1O9h7i82vS+e1Gh9Aw8WKSk7l
qExim1WznH41V29w59E4Payzyg4tdxLthMguZG6Hg6AjIgsBmYhLvwptG/aI3rRAyNWCGfXPO8sX
IHy9pOFgGXIINLQ5AkoRtOACsidlmHhPG+4u3kq11QjMR+PgJCL2KzVN0cwUWpeUPnWKdsUzx3hF
XPUaRUdi5kDs+zkyecpICwUZ7jodAqV+qVULzJdWGJ0cRto7M/7epa3AjxLoMA4wSKK1VhBD7CS7
qO+kA94ZJndTzRK5slup81QYavwShEjWp7Rkj9to90+sYae7fkTBhx/5y5aiEOHltmpczBRX7Yba
jo6tdOszRGR428ugBCbhIGhHQjLb1+WLsfCL9siYCXUNyxJHJXofLX2lEwXeQZvVODS86YWBgnTH
EfAhlNjc6g1TklA/bG5d6gsXoW9SwCmg73/eLhxMmWdP7AZmczoS+GHHBp+MGvLdDbCl+RNpTlSh
Sp28q6wuhGjpTTs7O5N4b0IR0Kw0xBM8mfmWb68wDrLYucbg8JQFmj2kbwlHVD8YXo6Wu41AcfY/
nP7XNDLZDlsWC/GrCeUj2pk6ZcH+lj+rXbENY3Xa/nnIC05DtwvI8Bu55TgPLelRfo46V56nKDGh
kCFX/tg+VMzaBDD5qpj+bJxBSGfh+3V5ltPTnstMXugUamhZKIOaTipJ2NMxPlCjpS3ohjNCgg0b
+jPJ/JqoEI8NJ6i0V6RlrmCL2yM35z9ey8SO+HLAP6QnVzzacAK763FSYslidOjhB+pSb0IrkH5G
mubx0A1KDv+kEUOfbq50U5b9ZmSKhTynA/Otm4zwXTtKOS3GnU9XSCOLWMMcHVGWsIUtQrb5vWqK
T/qoyAkdTJD0L1J1le12sQkjv1gC8E00hal8SJgUhWF5mRfp2+GsSkx0feBqYDFbtnVdn0PDSzY+
OWkVeOhk09vfrWsi4GIy0Br6xlnGz9F2R1psCkY18mGDIzZz22RdAvktJSBWYhjMYqrJcW/uiTDN
tiKlXm68ZdHKKGwW5qtxd+mqeIA4TyAScA8+bRXbZjavGebnhuASIyBz9zGw5cAemYfMr97O0SwN
wlxfS4K/mWAxCvhZdgQt5uNuIhHv4UVBKcLGx/3yvy40po2YFPc0HnPmBsDtn5q2LeJERufTmm/O
fXj5hHETCWDkaaCMLfpEwQsjy1KASNFN8mFf4+Hp05sitaGwQg1OE2BxuDHA3PrxUHCltJ4li2YW
Yze3fMVAL7rvfmZtkkXNW5gNWmhe6REJhmkc7wMYnNCZ0tZyQBD/cLo5DQL85dM95aqZ3mTdFzy3
4bmsRDb+zCjNqtCa0WaJO6Reuup8RIOKUlQaU70JIAZclro062xjsnbli5vgZuu6a8RQqj8cFmRm
N7/7wnLV1xFN2oBts+UlS3Jd5dUHPcbO756gPMLABFRLzLKUchKJPeudD2GG0lqel+/MedflpQSi
FJbPTU3Bpm86MLOKggMOfIGDzbbBOofPqnDXTMUmYQtBm5i7nfrIaS4N5aYJ+OFC2XlB1vX5Aidn
7Xoxt94q5/16rsmDTmVs1IMfOpGwuDrR0ceV1CRkIsyFRKPbJVmOJ8qOidiVxau00HvlukrCp2E7
ekGmU8vLxUVex3cIASWnj5St0imZUVe/Un+HnL1Qy5PZnX1PxBaJChCPJjvMER4mLpaZKrvXjefL
wqKpoQ7WnZ8pO72RCL20k7qRw3rZpDnmxoCZi1DIfQ2RQCr6sc2V8kDQf7DmrmD+F83HahqP7ChT
H0wN8q/i6EKsnkK+ajk1zEHZAcK35XeRBkvrCiubBO0Lo/7PP3YjmONLCt9aff3aVFeSZaXurBGF
8EDuAl8HHowqJPTm2ZedB/dQ2luYadO0b+RjLOCtEoyMbxtcZ69d8cSJYPGA5XgqoELvsVBfnKlB
fx2ZP4laFlzDgoNEMQHrfqClkIxi7O59gcCjsjDnRHXVWVnMWcywdFbeRQv1GGwhxGBhITMIf4QP
4KWkZ3e8rq/AU4TtRNRW2Ut/bi0GZ39Xfc12OP0ItP3zktZbRoF3vpzTW+bcdp1yIFOjMZID3h5Q
Lga6gS+HvdGgQeL5ScrfoggNVH8MboZhIpCqTj8pFm9petZUEr8E1xFX42Xf3E6LTIY/j0lFIrPG
pg69OrBSXkJrHpgow1l5oxs/sDl80CAs6PS6CKOiqqkZ0/D9hUfwv2+63BiADCS9J528m9aDCKQl
rASRTq/Y2UG4d+Bj8yDDriPIFeCKeigngfagj1vBlJWEslEQGkdkGfyJ0ORk7nE1/Z90pqvMdxWk
l6+74tFmZr/Ufma3866b7A8eeDyypGX8SFF4snem0zWUHxFp5bkn/7RbqsAy22z2QKGtx+dV3Zs+
smQxGE02QO8dyF32R+UpwP/4HspEpTq4eJ7bNvv2rkrkljMDhd4zIQHyWoMFb35J2lzxbAtqVirr
URqfAsCqd5NvOn0tQJmaqQIWy+rUNX8IWGafNaVSjSuLsxNCuQXgSVz9hBB6WQ3kXXs6kKvspmdl
Dl80U6MLtJ2owyJyv8RffDCXBEikD24LaC1DYuBFERcmLl3FLy+Z4YamN3EyPOx+Dx+wGz1xMeNA
pr5nQ4tprjxcjAIAF9g9/WtM3rSXs/lVWGA3OEtqiAAww4bJwMKuj6zTl2bvOTC1sc7xrzJ6BIB6
u1l1tRaEu9PSLguvCUcD63cpnjcfFF9oL3BeB6f0GjuLLjl+fxRXZ2QxgkfnglGvYVP2lJimJebx
kLtFQzh2n5F3P4Ffg9msllpl0xd4XtWfujMGCxa7tumFS7jT61s6CS4SqPvLWCAkJ936NBQIecqh
C3YO5dOa8UKmYgYl9jAi3k3eTSYlJxQD6OgYOTSRy3+LD5jhqRZ1pNlP4iOLd9zTcsTvls4afvV6
ImYR4UmnJrR1TT8J/hQkK8hbh3THsY6tm0lFNEyGQV4Zyls6yAPcbrojYaqccuRpeuUZvBsFQ1q0
zju7R3DtlyJ7mngjB2xgA1/WlZxh/xqdek1DucfY3IJ6Zm24E6AsjSZk0oWNIYITzfJjwFP4+ci9
SBQWEF5k/vwmsafoWETC5BqFg1LTySh/C1WLHrv6XtBEP15UNCqrcrDNt34jpLq1nkpgJplXtYTC
v8d6tTjLwe04YnM3vtwvd9u+I720NcncND88Up9k5GmJbWwAl5feO7MpEp9vgn9cBhO60Ej5U1qU
XNBrajyIKc72KiC0hcjUjMQXKpb4ARFxTknctDHpAE50K3ei1ycN0QpnYsBxRAIPFAZbGniI3Ws6
+s6xjsYB/7OPBOig589HB4RVCbQHHUwckPv0OqRWrN7n5yTLN2SHr6KxD5A98rT5Ioclgl/oqSYx
sPwtbAzL1dbECxwhtWK6yoUWZJjm08fAZOU5AuqWOoA543uzN7YPfieIy7ytEXdd//l7zD7aUZ3X
cCJZ5I/5JSn8qKjCLQDnUQ+ULJMnfpD2XDSimGXvL3Ts2xXoxiHhGGrSduTF/Onyx0XQXwSsy9Z1
FZIkufc1p/DA/aKSg/ngJ6flzSrKeYdVe6CDhEpm8qZbK9AueNXSRFBih+PxzlHMlVyijg+oeAg7
F0omqjBafcPpIwX8dfifWiEGbAqACadP3sw1IwbVPzR+UOjgwfYVNWwtiv8YkudyoGMUmWWUMQbl
S2VzArdmrCYF24Who62OAx7QHDX10+6rjEJSZ5EPjg4n8D1UwhJKSh3rdAw1vHKBDpjYWnapoXmh
fzO8kLMMrYdtlNUFECYelhWVHivRZl+3DehmGvXK3EXpHtND/dwkmlOI7XZk2Uc2KHnyP8Adeksi
6rF8W+gqvWgOe4NlH/kRbFYiCI0zSpEP2OJLLS9Q3DAE24CtdGlqAYy2GCdG+FzSFqAZSJpFvWg4
oSE4j0I2oEElYNz/Lla/B4OrkjMMfp6jI+294ophExaYfo/kfRV+QYikmln/9anRUP25JbW41T4Y
PMxL4S+vRclqxxeFe6eeflGfV+5Fm2t7WNwXYMvsUeo9o4ndoFt5qyqyeeNk947i5fKZSPH98Ptw
cV27UqTGsNlJBPLXdGlTj1hzqisoLdI7FTjD5Wya+Lqr0xXu4SHNFHUAx4bYvksm1Sujg4987FN2
qD6X7wy1BH0+k1jtIGV++8GXB+7BOLkoIOTsWQfXvVcdUDpXGqn+DV+fgmwnfMqzSL32YWJoQ/uJ
1DjJg3j14tc3HPj3GGOSCKNyX0jUMXQVvO24W4fu4pphuKX+aUbyh0JY/9gVXODRbvWxEyWoHmCN
sdj//ecUKb6jkx5PeeGpHgLVIFdx3HzOeHCFiYI4Np7u0qAMfhEmEyJwiqOJaEbRghkQfLlPNMBY
1XTPOA/lUk/KB+wkGE7/e38Dhv0B1kfVy83+IKIWduOyAWm9NNMU5/+RdaM2Y8ZQl5cykQGON+Wj
pMcGY4vumZ1IByI7aobXPRSLauEz8FPj3x4ELKQm4L3kIFpcMXwaaoRSUsu/qqQUFlHX+9AQfnjH
vE8VcuosJDT1JjJ8r4Vsux+hBSCatXbUvUZHij/eNCs+OAoyTn63GNaLQyhPxJJe3HyB46khUoE1
jkbAlXqEvr2dLOIkDC2GLlIZwXIpDIs1gzak3fE4R41b9WtUoDR7a7JDIvysZz0XwK7b7JSHaMlL
sSc9k4U/6uYoEwr0TvBczTQ1FuWuSiOok5VNGtgvcU8BeAiaQX2ZQfPTMbwy/NdTdky/b0oTPOgA
cTNvpVIUyu3T+4U8Q3Zv7yac4SrG9THQlcxTFm/cxaZgfCE40Aae/ae5wMQWWiwn6xo3yZar48Kt
k8vsVFt3y0/HNsUz9omKM5fd2h8ZOvAhdd2dExMtxy8tGdHl+Pgstt3GFck9LMKsylHu6V0v+zJU
fAYQvLY+3/4eUwx48M+4htzOPq89BvnMxEJD+y+e7/QiwhvGKWLelFSsOYlkyNWEaIX94VrzjC6B
4nVHi2Q3ZDOf+TKzdtH5EIZvHH7KsSUPepm8e5SFS4qQJnmjGpp/WlD5gFsBPpcQbP7Wx6ULORH+
JSTizXuFKYXNqZP/DMyJdWWUvez4EdTrHmSBYw/anhmSfULt4fgB1sWNTXHo5kckrdMNVt4w8qQO
jnKIdIeIA9JBeegqxdb9ovbU5Vwi6Mg8xh09CwL8OFr37shKOzbVQqidoaCXNIuoFiN911vsgije
do/8bWAqbICnRc1iMmF+3diGM9xSrhghRIjgEQaqTvQrgL26zNqGT1TTHdP+19Ip3Bz5YuHjr78s
F6Hp7sp0o1sLIAdtWii4b1Ddlm9w8vE6NMLcK36OUpERDumTAVi+9JfFrDDa02QUVIcibHXQzIxl
LVTZbaDj/VEl8yNAz36IYFpbnUgoQ968uupUM2hirEjpXw5yFTPLRyvhv2tHVf1X+Foaeva1e1PQ
dMomQPKt6G4DdULBKoDDT2bXM4n+fUDdTwKrGTqHGFFQAe1Y3kd7zEz4+GPgE+5Je05L6EKboZMi
VFYvUbRKTMVIdy8DADaYWdd56ylpMRiR1vxkCUmwGOfE2UxFtgg3BaVAn86IjAmCTsHVlYLL6aHv
EXFQHlvmxB9cIYRHzPK9mq1VcxZniP+/9XXBMnPyduqkJ4UcYZUPDvSXfx62UNhWrx+kNsd5NySV
va4AnT7bjmW8f0xioA/NCI/vU5+nvtYCwjsi0TNWMHFDBO9BHEek7b1PX59WJVSZ5Ro1CqRMnP/R
8gmbTv2GDcpf9t4yRirXnRkvbq2lCYbdezCIeO3N17NXnWghpZSxqsjKYYKzVung6EsoKizkLtO3
R+r+P1awsAWWHfAyppozdKSpHQHEMDtR1rWO2KyxNBwUMvSoU+ayEtXqGO4f5NjGizh6ZTjcnx20
0ANIhgwX8Xq19Dap0wIUeJ/6I9k8B832wviFcBjgigUfqa5HZUlxMH1/WLDfBFxVRZEEVwuDMEM5
wm8PAprwADXmrXhBGUxZFPPaarXXxgZJRkApKTn9oQkemLxSPFDpgjCypE/S5G8//+24fZ1xb4Wp
iGCs6pgqYvVJsNwtyx3g8+9Wy92z7NxWhLr+xx++6isWEc18cPL8fxI65dQ6F90zMvIuzVMMqxWO
aU+K8FKpTqZhLxcz2m21KO79SE/P1HZWyChYQFXCZNLcKJSxjhEq/lekeGcIvGA0mQC6DoAMgRV3
xdzqWRfE0NfyAVQMj5Q8hBKN/2PcoKFqVxFYf3ZvzRg7uKFkXL1wdVpMo+NOjIimqC4OPN+cCrF2
0qJtetwX2qGAE78VGDSXMuNBMrVreybizOz0aHQ++a45q2p/oDDOvlJv3/Sft4S64may82vd0KOB
tg+07MzPo18Y/FuzhlCtfeBcRMQOGXkAxeMDr4x/IJUuRn5luBL7bfWhX+LHQPckCpMF3amjll5b
tQLxoGiWzzAnBCWSCxvnx+n9+mRB1L0hH0etymb7X2GGQCV4WbGCoCLRhj4Z428wMDhk/d+QNhEc
a3rEofirNCxI4L14A4EaJUINoav8QtqzhsqNnXcCVuZw1afOjLw7wlor/GapQqSLVrCcEDrd/51P
hvnMqZD566D6UXmm8biCVmACGbXYgclW5onLkU8RckbqiQHR3tUZ4sQL5SF1unaJ1CQSt1qef3ik
sVQp5PJDHeFt3DZiVE5LNt53mE7LNmJ/gGb84UWDcxG7MPAMbYbNn20vsMTOA118OcRWBOJZC8ea
BaYmW5iU5j3G7/LEU4zDE4DzjnTkbx70eUSsIgJACczmxZtc5AiDxUCMwTMkvEMFXG+BYp1/dGtz
R8smQ8zh54RqTBzkL3b3vo7sPi+DinSHXcfn8GTtiVZOMsCFTBJlutg4l1Ng6E13r1uApG6lQjUH
TrQbqkow8MqqU18AW4trGqSlU07Jgx5v/iufL2zGAzbF7omDemeDhgVbpntxrpdzI/gFCxhsYua+
SRUkDyeJYdsWfwhsBV4DtcPjnIQskeACsTs4qy52Lp6heORYEKJ5lVv2ldIfoYlF0IOkwEOZSmwf
5540zBz4nlyFaA7qHThWijxKUx+Lnz/wOuLbDYxe3WfbCBJd+FXoylI42Gtj4UkA8zKJyfqDv+7s
QwKdrX4WLOX/1X12mh2g2jRkXb6hjeXBSffixoMSMbB0Ha2AbmX11vVx8BCPnebsWke792tZLBzd
QAxsQo1975RM/Fxkc9iFPBY51fb3geheNQBLR+ZpXS9aJpyiq7ZMcoZmtOqpXiT96cvYJS6lpObp
5HVmQ7L3BxZiA8W3PTcGRF4MkTg9kOTcp96ahPXYrlycDyoq639IHhQkbIANaHM9u01hHa8qRj7R
u8VkrEV/wpqe+/G550tTwxoP1HvBfl6kGczYr5XUO3o5FbYxtctlIhpwD9BaywDUquldSIrfCiNS
qaxg5bzAgHDYSdfz/cFSjNF11HzhTdJCndbHGlXbYZCQwaoNt3QTMMKpkDWxKru1euLfx45WMQOD
raXjzVwCSCTEcEegyV5FEVFTFdRd/tSw5G8CT5jC+aAY45C2c+MZczNLxYSPm8+tYdbuoIzlESUb
W0d9EYYO5Z2OHF1KF49wn4rNlk4q6imyuSMWdrScTTA6/3zPWD1A7SUsoer+6/ukt05KX/I93/Gm
pNDQj3FFndXpwMTgnLlFdlI/L3MJfdYntZVymNKQ8v+1LKFqgiDlnD2xy+ezCd20O4Gi836RhclW
WtzVBwYTgQYyyTBU3Lui4eSMh6g+EYNFfVVYKHQRxSKzd17ZqpzSjJd59NEVHrThNxBE+5abtFMG
9b0uDLJSrGd9X12ovYpgLgL+x5zy4/HDhbMYXk72Uwc0NJ08SPnJMVNb1dSG4xWDpK12hEISY9ev
ERB/mQeyatOEc+JrUZky9GZfND3t/HYGb+Kon5Kq3dM8AeIPFf+2RStDvGfQGV/c6bMFRbFuRRLx
gOehdRH74jRjMQmO9RoiyMcASvYft48nVIwL+Gzd6gE2zZWK++uucwjsVYw6Z26z3jBkIKGaLNpU
mdwY4ko4jAqjHEFKHAPx6WoH3LsXLEBDy+mwJcUCKWCe4ac1yABR5BBLoUKMVlJ3zBv5Gaylo9Of
EQaV82p6dAqomB7vxB9NeoD8fGoKhAP3fP6ecdCS/NcPlQIscLzljfsHYPdtrLXmz6JYkEEDWvzO
ghVjWcA4zsR9mJoUEcokAhqepIyvWiGCKjSqBwt8U33f5mQ4CebEBhVBxv1o+SY5NZ6fvuhTUxHF
fXgsUIhU6PDj5uuxsE/2OaDMa5Tnc7h27hOzdv/Rc/bppyvTXcIH5v6zwOQMzHqrzDJPkyu9D3vl
emzUGOJq1yuAcKMU9AmqEM1dOdu493iWA5JuLypErIBJ23CkcB7Aa/p8ElHIqTG5RYtr+JTQhQkO
JraUwQ4aIkudtQnDiHIkufTTEkwdlksZYhcJtQk4qMTD7SggcdtvPYHxsrsftYxnnq9WcRbDfhbm
SBw48pEgZOucTxaJRUqkcf4FtKhZ1ZJZnaQF2JC3qLEhWpZh0GarSiD/g7j6m/Ns9107ebQvAAte
k3OEc5aIJLYltTaNvsGUpHDFySX72nhpYqa6uw512zChOlhpu73LiJMrd/JT8aHZHBhxPU10lpns
n7d07Ogg64zIPz0giGWe9tGoAUXHs8OXV9LrdwfeFZBy1ORyFdOBQM+FOjAhPbhQ4F0r+Z+mXp6n
lSYaZOKRBA7p43TzcKiLhj/SUIdKapdAcah8RA/ktxffDHSmAe2slAuYk1dPV8hfDfEYFU7vgZDP
T8rW4L0VlTvaNtS06y0LDolN64N9/OdnizEmrVhRoYCP9FpKHQ3kyALcHG6IXNyZaEPJJ4v7/3WW
kzQub7t99NWMM3HZQ4UnbBUNEk6I8lhYkomTr5Om6foV+jfYUgLzyYW+FpA3CcOmF0s6ZdYRsydy
/lVAerS3ZuqU0rEMso2tuZeWPRwMsc+r/2XK4xKPu1qGhS0tLugfPpJR8dINv3zJXHRYsmXgdiD5
Hz8PGLOP6lOeQT+k1XqZJ/+eJR0uHAp05f9I5JqDaEVm3iSetArc8MfOnHUxGzW36fAiA2rLYhAy
U1tLYbRXE0Q/FjkRnL0qIowv1BP82dz4Af9Fan7LKAEj8CD3DCdU6v3MrpVaGP2FLaO6377ObW1K
UjAuNFqfqe2Xem7C/y9HG9D3HhhoJsdMFUgINNqxPafzu39BqpVvikDJ/rSxfW2luAIfjV7IBOd+
Nzn9/CRnUu1hnX6z599jFhm11Xf9XEUYoNr8i04G+FoHKp66P0PudMVWLa9cz6h6nhbkPCOq/XGk
yGsXaeghq9caf1fOEcnwvd4PLLP99jfj/z0qfsji/uiYu37L0oTE9+28O0FGQReZO845rPuZEwg7
hr8ihAPibDYSevK5BxKE/ldf4OUkh9lfc0IC7XvNhPTT/yLT/ogA8h8eq4+vyZUtFQ3fKNLlCTp0
g0TlzHU4s2tcuTeXYpQikp1Lcx/I85zg5Sl2UqsW70EvZfYMYgN2KuLOEtqwETYBVFlOwoPc2DLX
jgsbRHKFa1DFIaE0b8miiokZfXQZiSxI6X8eQnu4VQW8PNWSSnZKaDQUH5/Do5wDoiWq7heNxOAx
dcG3UNjrvChreUg6JwuRyCp3lluPVpv1FcMD/Ya1bbMCD8LZW76xet9lp8LDwGWmLRMhyWFOWaDx
vWeoKcbfsBfqZnrLcS5ibPTxerbKaJY6RoAgatRdrb5SA+ls8J0bN2Q3JXr0od7X7Tuz7+6QQa5k
K0VssfJgAG4EyN2pTS5S7tftHXaYXXhL9TN5aPCPewtJOC8D8rM8k9+xTI2xRIeu2pznUqtjY+bT
KV4UJr9EhNc+5P2itmdmZAfHMWf9qZ+IeuUcuiVAcleMSpSae74NC7co9cMAay7IiIoeWm7vpQvp
sTEgyVkvOSrbOtE7oQJIL/ISFfo4dE+XMu+wBbEQ2Werp6Id37nQr8nsUpCLEWK/wKyo5S61CJzp
vPtj1zoUzioH8TMvcYm1/+/uUXPKb4v83j9f+qPHSmnWzaoNp2YgehJLlRL+ice788cVv4E2Ynck
HmYwEN4TosdKCVALFaUQyfL9GOW6SvWPL/9bFcUkXaYrhAsR2Y4/3eaM8JtSj8D8dZxno5hnDup0
bArp+nDMpfXyjcI1Xt95t1rVhM6e0UV0I2GEgM/FxyJcqniFupXSee4Sp+9Xj9p2UWJfhoIWqXM5
zrKAVLJb4pHLmwfKXWw407ryS8lXcmHS47oWRe5OUE5XQX+YSF5taV/hVBS5rZdcNgfpuDBX9IJS
7yHLsq4TNuxj6fEcXyTwsjRLPBdmoLG0Hww6q1AbvDtQM9bAMtCFXQaOwxkI3AWLuS5zS25Nndm/
+JjQOwQ/xkad1NqtiWelXu4CfZ7sXqf0HbE6jkFL0sVjzOw9javM1j0aQtgvFNTEaPVnQ2GQ4ZrX
sj+Pz+oX5CDphfEm4YDgrVG0dtCFdbLDxRN66Qz34l49o8p+9mgUxTHoKvtsO/+b1nN/IqZjkLL5
4tN33jw7bzjHmRlp9WZR2r81bIHHLV+Nbble+vqx4P9FjjCAZevcrI/bt6ZSyoUSiiGzXi9TG3hQ
vAJE0GWXBlYyPCqq24PphYx5BQlOUAlHMPC1NBPXAd+rOH824xxPbANA7uBgJPR3Uek4J6w20yrF
dJggC6H9ZVWiWXbXu00ln88Q3qifETgX9R16U8V8+IpSy2vC3Z9LIsSYhEpnj4HooAVwHPIsO4DE
WSj8JkDWX3IWXR2nzg5kal+/10EEf+J/OEgjEkA1CFP6Y6WWwTWq83UlsqoEXw1E4wOjuEqDvj0P
6Ai0PWO9H4i3gM0R7sygoP7jnnOrMnt9bwOJ1cGxUzVHaBNo29Ee9SkypHiCLvmDk7VrmSi5efcH
HC6GqNHvTyQOhm8cSl471Rp7+a45quWLod0gLKqBRbClsww53ecVz05Du8tQbWjRmnmWOofw+OCU
twnKoiqm33LJdoFJLFZK4bCzhbAxPmeqtbC862pBPX2PePFmIOEqZOftZqOXqdKhLeoAtiig4c81
KJXs8gwYLfdt7E3E+v8WBt3qkofyQyMQtDzf7rKc0EDLde0a3X0eH7e6xuhx+sBqMow1VB6DlZsW
6mUdp1C/qAeLH7hNgqjYjlmMcsrWjKnIbF+4won0bYE8zgHN3fx17r6eKB1gHZU4ueIhBmTYonj/
sebdwgPaVMEaM3PabyHnzc+mf9MivdrpOLcXnl+p0cnyee6wAaab9Hg8jnZJPgZXiyjG/uLgfocD
bNfyeUyJmwNVg3YZGBp2gIeYBpZsx4zV5P0+9NByAbNR2JQvn1qbBjgsRAJ6OOuvmQGzsn9Os7wL
QX3aRqzEmHKHj6e/DC0cKRYB5+Pbpnuko0+a2DGxuW/zbZiVsa36S9PW4523sMZRNRju3CSiHRDF
rvFJyNsoqMaqxVVSdMBkSYC071117LB3prW5w8Mk9ZI8jl1eDazCYt9xXeaAg3ztoWEfXOa3ML81
mGmFF1hNYNcCwQ+ylTqBzjZbjgCDirP6DEeBfaBpDnHB4ys4Z5OkJFmtYJ4ZUC2miwhE2jF0oG+v
SorWH2ZV+/F9ZYJEDPHFWsXvLe+fm2FRalBTd101TcX73HeawCpepnea86chsfYC6RpSG7CrGA/L
fJlwTNMAsFjt68QQ1D0AXSmoY/IfMCPrP9h0vaOcdkwkCcvLSDV9BZcTYZbb+HDcRs8JSv435QId
N75k3C+zxkbtNOjxKECrnQBTf08QqxtSKmQFccP+kkDlwBnQeYC8XJ68QTVoE2oXxwVSwY3HX/gL
x6lbIGk4LEhc+CpBHEy1WijuHhySyq32i5MG40sOFFukRwKP7QG01sAgzu9LkIGnpYmWnzlRxdwQ
ReCtP/4dOgkhm6NnW1Y0IMf6hip4gqeGr1ti6b5MeWtdkXknby/p7JyB21xYAxRqKDDaJnBP2hMs
mFJWzBFQxHhBrcptRgBX4uy7i8uR9cCQ1rr8Bx/RXzVObcr3yUtLWQARUTo6BvGwTdyv3YGL5Ge+
4QU8BNXE1QU/+O4rw0AKRoCrME33mCuRkGemkCEpX26WsYT9M0yVJqLCz64eQ16tARrqmFt+OIz8
dAt4YKi/aoPYLi9cXv92omAX54f8Uu4qSe13fnqZqD8cWxaT69JaLOgCRutCG8TBK6C9LUbvXJTw
IpbRDTUQGYK/Y/TjH8dKBJv9AzHspvx6QRfnt0OPJJ5Hyfr4pyTAfupPzihQsFt6KiRWg3A81ryL
LNXEpnt0tpRTgN36m3n4UXpLN1LbmNHQ7KkFuF/l/7pZE2vt7CNGJjdHiyb7kaxXoO4aXVNutHEt
709Ic260HJ11hr+V7QZ7aCL8mEmrPIhKtn8L8szZs0K9tTASrVWjhPqHk1vRBHjcF/E4ak9P2WZV
+uIBrb8/8Eb2gdJxjLEAMER+joGz5d/p3h8gqOm5vdCVxwpPFQLt6secRj2p21yJeeV7FyMipie0
ULxDg+/Xxpnw+R+UedbUTfky8a7bnNTCGj7UWnRlnRDeTMjkWuDVtX/jaHyTcY6z0WHHKxrCYubn
Ub50Se/NVLrFo03671iRctqCwWPlb8UJJPNOkb0FtDVhjFAHzuD63RoRNKmlQ/xj6H6pkPyDDjCq
nbcr3urFpqtDvtjyDdX9xvgRO+TFJXlyTUX+DDrzl9x73/ZXBJccLumTX5i3IgSfQkwNBXURSh2H
hYBNeZZQJY5124usNAET7ywmyOyd6S1dW3sTTMy8jseyyocPAUr5lvqY6y4Cp/vFH+SGXdG3ed/h
4NWXR0mS2EUMNoQGOCtwR8wumyywVFMQbbp0s31GCJwZbMoQ6Us/2tRSqQ9C6OiVwySYZyhzpIpg
kE31CPJSb3+U9qdZgYsgu9LHGCzzp3Xj+4KKXgoah+Wy6ol7O3Mg7csJkXJshXbIlyclZfuIiBuX
IBP5gCKZcgsDQjMUJ/hQWQ2Fa9U+cek7OzEPn00Ng5FMBF7eH+gfflZ2tSOjnqaW/dpfrZqVczuG
3zJ9rviWdnU88t9ljW6mjqHcWE91JLXdZ9SFs2AMKu0qCJQOOECxO7yqyTHJUj3slwm8/fOQ2jWV
+b2isL/lf/LyZlrVh3ve8hiNpvybUSsC4aKENHkFZZxriCy9eHQCmeuZExjPwelBqFY2dy/2CYHO
Hu4z6X62oHpul7dSYt2iNIW2kJwCWvSSfMxw5SeQd6JTSmlVOasXqfHhsbZtB4EbScesyIGvYfsc
TJ3J6dSglBi8jpFAR50z0PRIFxuY5pGshhP2vscwzbieEpswEIcmb0CA+5G5326IKHj1JQzplddp
NlKQqfx8GWfUeTFVDRc7GQiKHk+j7tWgWM92MpChRmzifLnI/zkmhtjxiRzx8Id9SMk9ymkvVzPK
2xUb34KPgDXM5C9DhsAOhXyLAzj9es8ZpLD9iaAPdQy1wRXmYpLLbttVorptsYRemk8XiH5MMGY8
FTCDqTxtvePCpkyzKFNd9FF9L1DURVhd2OTVtBIUJKXpNjA0enx8rULGwiic1EL3LxVk8NWww8ft
iu3DpS5R4SEDK9u41C5OSt7aZs+8PX0RRW2Ad5WQ/5yV6KJN83OTONYk2DKQG8fSkGcWLEAm36bs
lmPO00H43XxQuSHXtbevepGqPB4dlmDRnc67HcSiUhTdKhX1snz63f2OqTVgYG8Do8u2HxqyfinJ
YDn6ZAeoAHajS6M/Xnbr8UzSFW16sBJzLmx7ZMNt9LknquGwpJX2L6vaP9g0jQhsatqLtrmGHTFj
fxYVm7+s9WS+xZk44nuFUaUTP/oqcA2x+6l1+OOGiKs137mS5r7U1+RpGSfR2Uy8WTlcWOxw2HRE
x05KFn8dgs5EX2F2zN09f2qtYavHez2QSWJgupNwgLCzqilSaSeSCpPi04bmiIUjHjaFn6BrwGIE
NBVAM8KZepOtuOfjqFaibDn0yoxbg8ayPCmoyXKKcsvjpQHLxIgrX4g+fYwHJUQO9bf+M0RtkF4a
N1DChFBt6ehShNKvnVE6ZAXtf6KDGFLxvs3WhkoJvy4Z4e7/Qk63oHnekAdaWANnmqgEZ8NAOVR3
VC5RoBcSTugoqPVil1zqMwid5wnatTzuY4iFpnAMQaE8+wJ/2ShQoAhlY+hwOk62M+MmTWAVErth
TVH8+AO01G2d+QFlWtjhw6njpw+Rw+1wq3d3QV+ub38RSsXRiVxzpDw7ezrob277vQDsPVPrg6dQ
6tiL6OhcxnL+XarXJZHFAsTVfEhDWlsg0asstKAZXX7AEuC2Sn8V2ka5qRKoOK0FGGvDe/Qd9QGF
yxXK24QJskTn7U73p2C3cAFK2qcU9U2xlErXAJRizlMGzjqaRXFrvsAFaQT43MGrYoKaHiQSW9Hg
VHAw0qrLfmyUMixP5JZJBzR7hkkjwy0yM9j1ZYbF8I22gWgAH/eccSDXHjWYYPxHN+Hld70Qd/go
5wT92CQ/bkkxj3dl1n2FF7+l704lWUwQ7pg5tMv57EXrqHuV0QFhxnCmNTLsGDBEAHNdb4wVGvYL
nVAQYIDgBCmseGCVlZpGAtUSZAL84kVGJkzRwKDw34HWTdD1uxc2K4uGfOGDwUvFT/FzYOR3ISG8
VUHabHquqASXDEvQomeHc+uNAYZzAolnSfc+GGCI8Nbrur9O2Lr0PwR2tCjpBn0tDgh0Guiy+k2+
soXNp/yGYRd+xTTEmEfPo20amvzuhnngRh3TE/NCAINSPA+MUaDN/6rcv3cY3jADSvIy9v1v5MoC
w3fr1fppsb8N9HVeM0Y810dRnTnUgmnb98ERK67b8rW9C1dBtHbeE+aRnBiZUX34VszWvS84SJW0
68iLWEiZfOb4E71h+Yk4+2v+lpk8LsAxm/WZwwQHHlgG25QEoSVnsUxU2d7lG0uRZRif0Jq3Bpev
PkXYbax69V/3g3Cf5kSIDI9zSmxkAp7ureBXTmf18L1laS2j/hRE+y6cvdDjIcysjXBDqzZnbt5d
6KPvMLTptbCqgi/neqhMvp+u32SE7hcHOIOS8gduoNe2zeJ0njAlbBBRvzh6yGLEULqreRIhVt5q
IZwhzp1NIxijMefrsEIoc2fSqdHiaUgHoOzrcBEIexidZwS5e1G8yJEs9Z9Pn05U2A7ae1cjQM2S
nFQ8zm1BRCX6+hzZN4oK2hiSHJzc6XJxh2GXhOs2YXQ1xJGNQGY/gAGC3X9eTCxl98QuYmuH//3H
LTPNKFrBz7w+jgdIm93Z8hVOdmAsShXrl4qzNVpMT2JnxDVH76pd2W/ptcWz/yi49afrl2lQZZY4
YvUrsczAjNdeXLS1IJ2ySKA3iYV3r98DyvB16oFNeVkdsr+8hIZtFt/xowFG3Y7Qp4n6HCL41UDK
ri685EVEBMNRP6ee1Vafrfj8GbbPOrOiJyH8Z1Ln6qVoTocgpllxKwDS5FZBtv8Szv1Bx5XuKwJb
YEx6agurf9Z3RDGm+TWb7PXVHlkYaSVMCI4QWuK3yupQAU7auhm3zDBtc0r/rG+z4g+z8t9uNvN1
YXmJM5HQEJGuIwH2WN21O6G+CY1D+l4kdQ3Cv5vVnETqN4jYsLQFw+av71tKPMVBS/jgcbm2MKjm
CWPoLVnUTtrbTlDoLtpZbuuCMtheeXvaC5/JYt2F0fVs9BBHYzJLqsHN9gu1ZUaF1lt1RQZjm/j2
HBqCsp5Hzo6530oIuIpefE2r/g7Ixe0yaxgdPD53Dw9yCJ4ykxB6G+bi+y7/Js0qpPyPN4g2ErnH
e2pvV6At/3IiKtJ3HZdBVT/NGnlvwmKHEAEcQSmx7CgpIU/RuLxVts1sbUcl/sV9hbYIlXkJNwOS
0p+RSn0cAwCF27n+2Jb237dVHE/RoRAagYfYO5meNI5pL45ydzb7W8U/vU0hlVVqfDSs8FEgionW
qvR1hNvlxCQoJOssHGM3WSRe6EDaPCIehsKUDWvhM/U3IYr4MnvwyjlnKk/LAW5MVB5mLpRoZPtx
GbzUo9klx4wjn4L1uuvoHXObLe/RSpXOfdgF+203JRdaZK1kkxO6r+VaxJsIK9adWe3DI5FpOycQ
z6SY39kbrzprxo7UBzcvKU500M79gcD5eKTpest4hja9xMUGdDo5t9/UnaSE6UUFR/5l4sUGh2Lp
3QZ393curOequ8JsJ0IjJ7qe/Vi3umGXi3FAw8FckOCQL16tbQKaBqGYQQ5gjBBlrSWk3WL/X2r3
pA1GKTryogUCD+RfAJ16XexparpmVL7erSguldXs10TEv7O9fwFVeWUXz/MFM48PLk3qpYWPWthy
pos3fz2G9m6Mw9IPjKHNr4Z3mDIDbBPN4Q+k/9UAIq1nPnddK86x+icv03BGgYyDzleVXr5QWIej
eAEN5ycfMN7zFfYP0ULryBwGSbr3C4Bb8DVuDdVEExLnuUZfC/Y+HnjVuL2doRkGHZtJunzjACaP
iNPKs7ofigZqDRW1MHxgwrvrgrLwl+au33WcPiySOj38NzEUHQSs2cO+OP2hxLMPaNbM+AIkjJnz
i5yaLHbyT+tz7F8zyKOF+QDSy/7DRwBk8Q+lM1Vu7bcHneG1EbGTukeAuYV3vaIXIEdeOhllDrac
JvykGQOoKW/0IUtn8J8JWltwY+uNnXQrztPcrxCkvgT+QtEVKsTdR1lY11O06r2rk+aW2+y15oU2
Kj1CoZJu21ItYalKBNn53CDMpLI4jW5jfmp+ij97LGXxNsUlXNwtTs2S1fDbfXuRQVFYowIuzZUJ
XUfEaBTXLB/uOB0Q+jPfaA5nUpG2JXGCwDyRLbuZgCRqxdb7Relhb70J5QHF95yl9kTkAc2Dw0UG
CAa1b6k3g3EVhlcPR4rqChEJIW0agT4fmD+r1J0wQ02WktJy/BJzsy3l67OO7/O5jzqraOni2zK9
s0k0PuMhV7W8Pk5fDNNKIyceFvjGTPFCuPwCwj1DZp/+j56yvFaqoz7ipz+9Umb+IuXlIDZreK6x
xvkoKnj9R0l7dCQvUw3DBaH+7T5N5ccO02sFdA0NykfMqn+EfSgu8DLFBYurfj+Z/oQ+2O69Jcn0
UMinb2xKd1wCm7Qv8v+eG7v9/+18rp3WGnQMD3yxIfCfNHX505Blbk6IbiliRs2THJahmbqs/S6v
ipCJTRJyGkrIZw8elfSoMiWv7oKgreOZshoYt4sx4u+OMdWrXyl+rzfF95lVcZhqIXPrFhH6C3Qx
tpx4EkUTuW6Uhrg4iyC0Hp8DQE3TUl+3yQrwDmAErwbSqPCMuwfkMR1aE6CmT32FXCPJonrSGwX6
EzOcb+dCZS1gkPvzPPs3t5vwiyNAs5vmRJDw+jocRRStO+/STuevMmRljKHxcqAHC2LLCYCdUIub
nzFp+oHHxL6G7hRlefcn7JKVs4iFUzO9cH43HTmyn867qqWKZJbvxeoFpki0oIaUFdW1j0BMG0pG
5MGwXy0WuJmTVOOveev5GBMyhlU+wlIyUQeqZMAGYMF9shVT75zy0T5wZ+pWApgiXKGKZhc0+L5g
ei71owBHbhMRZj/SRpmLDA6RnyfG81HLBukmjsDangdJIORrvD2O2nK6VI7FJ6Ci4hVDBn9xqkdf
snMEo+E9bZ3sPFGfuQUlYx263esq5nTboylFav08D92jVAMjN2WM7WEMAWQC2ITWg7nWgttKbHHA
hrinS+ET+mWf2cN/Xn3Bg+KrbSGkNTM+wIL+5+0w4Y2IeOTmx94jhIWphWsOEDy48R2cNl7DnyH9
geBwSqYI8tp0lvYpu5lGkOIl0ezk80w6FkBbcwDmJizur/TdYmjKcnCOgfyC4GYwboYta1rnL54q
OxtLpaVq6uwGcWEAWzhQgjOk5uleZGEWMmqyZPWAXKRfIz+Gxv2X0xreByyPgc0hXz/BS4TS5jQQ
X7c5SciXjQh7/Jw7uvvc//+83jwLnyqcCg89hyhDJo5hQZbbYfvdjNViXw5GmEoM7hrPlwRfwaEO
l2bxL+QMTJDn9KURbyNQjhxoLYiA071IlCsrZJ2ferL7hK6G79MEw0ZmBaeGv9t11wF+UWfGxd3I
YjSUwMAFAmvvv0SsRsBxWcNkJi0YGg/iZ2JVH3HdWqI9T8VHSYx/XjIlWfBejORUEGY3lMAiTOWr
IbwsHpRnXk6fe0YRNMAWyK4eEwtF68CEDlxXUfCc9Wp5BZAalJta2DDwCTD+fdPfMgcH5vnqVv6M
HJO0rvxO7dFFD7d4cXtTXANOj5UsvFWAhF40FDwVLROUy2wRD1mc1kaF+zc6cy1bKwKkB5u6yjhj
rsOFnbW0zSomuxMB7m1KfDNZ+NTbqF4eaL74xn+nij9V8948I6mARW+2ONdmPbfmLBpnrwx9/8hF
WBHchAZ4hJkscr9cyqx4xPmbglBeocarA/n6Bur/j9LX+IJn967qcPoWkq6+fhuw1ZaXFRjQXsIZ
PRHxAk3gnOlLvh6bJ+YSLb4zBNie8fTvuEDXf4iGbL28qfZOl/xu2JXmtZhj4Dxui3Ne+Ickse4y
NrBl15zG9LDLU9Kf+kWFnjDXK8R4khPvZsaF01uutd3SgQWc44zNoziI9kPgpDMf0NRKKYj+QJgY
9r9DQAHDim4gbEXHIclORgjWOdHQqn8pCJIF3ODmwI3QKFZxsLStPeKu64fDDu+kJ0NCz76Oettj
O1f6Lh4tw7+yY3kMfoCwiE6FWKD2mzIYI9US8N5SSuy4kDElfgf0p7GC7uG83KoZfpL3dbK44wyF
0ZnaBsVbMTO/oxiqavZ1EZnBuA7HyOuhE2Y/RQgWShZeCWhoFpZYXlyONR2flCMog0PHRL1ZWDFL
B6/AzdNOT1Ilpo8pFwLVP+74NGxakCJpygI21Qp/9WoAZexPA6huSTb5Djl84N3aRN1NSPvinTmy
q3ftOoeIfjsyML3mq0uoIhshthlk8HK8k+VRobgXLKPMrk0ruS9gqVc5RFHr67BxEMVun2lX9olr
dEIypn+9UjG5dWtmbcGkDBgjKkjREz5FVqDK+vxydvQVzfFHIyajCEPcxncWd+Wkv1uFnK/QuV/2
x0o9Kd8uC4gfQ0c5lMDoB+GuFQZI7Y2Q+hHqfjeE/2R86tmQZHsOQTemuKyv6UAVjrmOnkXV1D/t
w6tmghKOEcVeaQcIY0ChufZJ+81d3oDzrTnkUmJKR/HQQdC0H7Dy86lf5b3mv++YOuBtIMZ0uRnC
yrPDFHsE27HLGrC/1CnfjPnil1KmNd4iI83m30nUgrrC1V0dfmgz0ivxyev4OR6rBLd/sk3zfL3I
2Ngpxqep0zB/FG4L3Pb1rbPlspwYEl1pHSkNH3VmNUqjK3j+AXqVSpWnJNFdnHBzNzy7R7wuPh35
m3HNOzuiZUmzKjt6GR67jWtaTGXFhEaM+uc/v89WoTHbEkaJgyjIyN4dAv2g0wEantUguP9WPkTr
RQVa+GLW+6eiYZvsvZGCwBkjCVuGpM/QAsh/DDHQ3u6/gw/MtPrjQ+VL6Wdmj3ahn45TsupN9mgR
eW7zXMXXm5c3yG1niySYlkmM1T7n9g+2sDwNy4Fdhb7a9Q6MZd0Ib5rfp8tI1gFe9ygZ/g5WSLZ+
NET914N7ocHfbThe6SHYk0DDhfoVMLAwhN85Y8gRPSw+lOacuxeUbMDxvm+cQvL53Yfh4HCv8MfE
RUPJ3hbiXHh6BHpcmjFc9BTAWMVRut6QY8rEg+Cr0eWOz6xzrqRvgTHAh28sl71rvRnyd3ZTg+AH
jLjn0bt1W1jXLTjoJGdGXFVOkA1tXLK4oXcvW3Z63jj88V2f9AeFB0KPvOHq5elLgXS7sW3hYB8M
aplET05QSFZCJvAIxCtDOt/V9SQw+Jr5o7IYC0b49shCekb52gdJqYxbItcDOb2IVSssVzfcz+N6
K+EBlyH8taH3LRb7EQBlM/R7w86DOkIz3E9QQ1aTq8XZJ4JIQUVD4LHOggT9MGqDkbyJoY3h7rNY
+y/roAEWCtN3OCLiK3INIXE0/Ros0Mknokb7x4nzPF7CDv1ptsDx/U977rQeLokxsM0+WB6HxyXR
Xf9y5yp5FPZ5EAYYhDBoF5xJTLa1wONqvRI9+eID9mQHKVzs0zd4gjwtIStMNiLDvNwrgNmqbIcw
ivPzuxxdW6ikuwUXjCeVV4838PjNHG0AhIQoZsTYH9lNF1kLJu2xkCih+Zp8j4+4ai5rmSsyp/Dt
AnKG6t8u/YYiOtRBKStLJpHEaaIkhaMinThVaEP5sQtQzqFSWzLeAf58u34QtQreKMA7ZnPIK/iz
elmn8fdcdmrLOkqasvPZdrKu6fRfCaN0lcpSUvnEoxt+3JhMJ/GBgZMtTUX9aVqYw6Yf2SoZuExM
xzwHACpsgRKwnGUf6jxlNp5n/LKxoolZUEfM5VPVj8c8pIBNWu0w8t6Jul1xQ3ZeT6/tYc8di9rT
4Rp2qrH8p3kAnG1Nqptn+rRX7A/cXdsMehyq4/pSdpLYcaM009Z4z7NuSXX/+/9rrr8tpSJ97/mH
seDMRtEAiV9bDsLPIQz0BCBNj6ehbL1RHCWhBEHjljZi8j63UUm+2ub1waK/efusE8vohswdifmf
QFXOyXNj+bzFJuBpr/KgjF5s+bIAu7ZrgVvUoxQXIgyUbkapvOWbTWdkWXz+XuZMv8JHuJ82udfs
aNMQdkYYkZRJznm849pLywPzV4f6L9gOCA3AT+OLrL2yZmfR0/WaqRHbKwBViZQmlZk+ehW4Xgvx
vGKN15SR4BCoT/R1futKKQ9SO/IhFua2ZugUCxXXi7G6JCRqsavNtaonbQtHAHx9BQ0DpYhb6ukG
useYRt8h2uBscAerdM27w0bnH6tB2WIwkOZY09r36ZLzF47Kd+js/qmqN4yPIDtkxianfdPIy12e
K2pCLKWduI6tzDXJRJS0jJ8Kb9J4Y22IGy3+jxvZvtBM6vST5gcXmHd7N8bxYRqwRiYhTOm91x6c
pUCt288G5RErzbg8DKu3hfNOjWBJMR6d0tUoPIaYBMKbxyPvoFFi4iLZ690xrTJgQMEh0aeojyWl
gZOqp0yyH7z+P+R63cES+qk2S86jyt5ARbX8nPSG5HFMrdQbr9lW4DKahm37npRR0SxWQV2VilIv
rPTfSoCzGDdjvk/NPF/UHVIkKGaLdWt9SAas1alzU1F23n0TNRIk9XTwpmZU4WuXdmiYCe+KG9il
+F9g2EP38i5JCZfs+cou1ghnTpEGdVW1pu60JD+Kz627NR7jW2nnwPqAq7KCf2PnCbhMcGniGOLd
55l/OqzNK8u1PfqvYUGfZbwcWFm8ujIx7U9ISRAX8nygZAmAOF9ajof3aMBnJ23ORJNRADWdUDMX
fg7VjoRafI3r19JJEUEg60TDeFo/cgD2K02X/6XRFmZhVixSQ0+8nmk6x0OnIqFpoi60y1UznCqm
Jv/HCNNOOBISS5EcXy1qptMTimpnMio+TLYED2QRRNeGVx5SuaAaknOeFvNsNyCyD4XeZ2W4oxzq
70qBW/0iNsHd1hxjgkD3IoQDJbeXjXRep/tYM1ixQ3RiGk64O2uCgl0/3XgCuhbwnuXKji3tG12v
eHIg/Jpopj5aDH4TNq0cziBfFq89YlL5vWlSJUKZUN+s46omMtGWk9k62DLe2QjiY9ZXOMyJg34V
nX+vtOnTp/57eeUJYFrf2p3xrhOnqrLXtEgUmqyzYre0kueCKQnTf8Bj4cXE4e92F4NsI1JSnhMM
rCCDm4oYWut/vB/OxqKS8UJGTGlpk+3YOPCgijOCFZK18fU9S8GjwKCbx3xSWeqJzhEGruIUjTGs
eM27UF86xZ03df8JuxqhS6XpNTn4fFOLlxC1JibC9ck1PDaMsw+v1hG50wzCetiQz6giXqoYkGES
r4gfaqCIHcBT1/CIvZhOzmddWsmfCoA78FtDQnDn/Au4YAJvM/L6Tgt5Teh0WzGg0TyKwH9hZMcu
/pH20FPXBdYbnIJygz8ah7fYi6SxjlV89EvAXusbD16kL75C2mCP/qu3Y+0pvXOnX3eQnL12KcWn
f+k+ziYGgcAqgmHqRonveH5dH4Rk1b+Ve3Ucx5bibSVsXBO2sovXZw6/0FuBCV367n5B5eWSOjc1
gk4TEe2jhe5q8/5c9bXUFyiHfQURVbureniqZK8nbfj2jM4y50/+mkaT29P1x35dIsPdPotglEaD
8kiJ49PZwwGnXfh3LO/HnDJZ6PDsN2FJhL4IcU6e5SxXTZ8qtxCdeIKnzqis2NXtrBX4RHp7CDHd
hWw1NrLJjWH2ZBmfUJZl5dWDv77zy51P/H4Zw7lqaNUvXadNbJ9BIALwnizgCkj2r5iuj6vNhg8u
QYiZJZDj2eQhCh9Trt50NZx7Pa2QXK0mqxKZQ7jemQ+rXWHVhH+5DrgHu3Bbz25wTkFYkR7c2kxh
awx8oCjJGp5qw6oiax3lXaE+BYaXrflmjbNQM2pworn8pEd4UmdCdcDyeMgOmaMEJmZUj7OpWCQ3
PJEDJao/zD6f/5pc7Q5Vq2DjZoqsEDdsHAtLE8CvmSMYHWVL/dY6sOwCMnYZK90AQETcrTb7T4Zz
y8tdf3z8HB8aMBVregP25AM9S/oKGnmnfDt1ROA+koBwoISO5sKVfdcW5GOahlwXEfnHSi65nVff
wBaq/qIA4Eu/1+LOXXDTjmiY9s5JYrNXVzJ7hmOWtYa6YkuimVDMZT7XyJpp2bs5a5ZxgW2dTQHV
7IeWSSx3q1oxwC9OT4TIwxPxihbY3qMyy0qCS+uNdo505YvsxRDALntyvc49Nq51Ri5QMVaJ92sB
iIq1vAv+WO9DWdSVALZjAg4XDFQ1PE1H8CHLr0+RjqoWJbQZlod6Xo2BfjqEAS4xvJWEQPZvVwgB
SSSG2icbxHfXn/YjAiVOVpUxgvOkIzW7AmRydB4SZg3KiyuKm4UtDPa/nBsseSvKPcRNepEjDt1q
4OzbWjsXzqFgGvIzz1VGscNlX6XUnC/Yu6ANZatXJzreSm00jYIIvzHDxSHpMLBfTmCffUxSg6mb
Hb550GmwfGtUcOJwtRZwWTP+YopTjeF9zkZhoDveDXz2V0/ss7xZ//OCuciKqIfZlZIsUdIVqdo+
y79/IAvubcXABcs9PVbNNT+Jq1q/LYmQMXhSz2e7ohUCFaBhN+vpQn4z/+iyPtCgvjRrA3cOuMZm
gCnJxUGeoXzRg1KcdR0C0MmU9XVswok/MHIRF6uxumLZ7h9SYR7+ghzqkxAjCC8SI6LCkY13ux+5
Oj2HQoKDOJWTb9y8WN69IBWGakbD6yppriXeQlZhMaXfaTcIwQ8s/bpo9vR8QcVrEVjeuesaUOk7
Jz6FPPVQ+GvoQbAmzXFVdDCsFcwDcotz2pue5UVgOSIUan5P/Bb5kMWGnBUZL5tdZrOfXTmarTjV
c54P3GXxow+ePHiE2lafbBUBsNn4kx+du+HLdy4kDlxbKZYgQzveTEqeyp+kc/GVqbQ6jj5eOPL+
yLqnpoctzZqLmDWyU+v9g5SBCSBxC6Tg5HJI45olG1n5uM0yrowZSykk8+aWTvySmboxMUsQSczq
AVe1vlCwIsgwvq0H1f+sRwwDziD/D5S3Xa9d25IU8wVx+5bUKSjPIq/Islx2tYt9TUQ0BAOz6lHH
3hL82C3AAjH57h/9ZOA1+cIV+7oQoIKJOiBAXTniAwJL/3obIkc3D90qO6CT/PgPJnZ5+bdlup5W
15SJVbSuBQFn4aX+b2UzFVt+Jvv39QM/nv7x32iAWCA8fH1479hiztWfG0ucVTZBOgybiwV7RH+R
089OtT/jGbZND2hoiI0NqZ5oe88AtcvGR9Rh7W1U14TtmUWbFDjnJu+kxMMusjJv39dbajDWGVjy
wTia9DGGcFZb9/ixn+ksZQZSuPvmOufoI0nseH/QC7Jtx+qmVAzauk35GU/OyM2qD3FqczB5tx3/
RW2W43vm0sZcm5QFyie1xjpNsdfVMoV6hlZr8mKgBqgtew4mJ7dEmla6LDAHsZJS5hzly8Vd3bvP
+7gio53ZOlNeGnA3Csf8y8hdbJUMpmYoxWT7fPdfeRPjaGTjgNSXCPbGRGRuTPIslqQRq0ir/Uvb
Sl7K/u4GzDCzZEbqH1rMaodjRJDr7Bsha07hXzn38v5z5yvEF42jw57QCH2GSvShkjdQcV2c6dXD
Dwfq2un+aW7ee4zzIN1We+AQ9oo/luNVtd9zI3tJDWnuGRUFKBq6ipCuoD4+Ktvu+Fm4H+5N0dTP
DrdFngrl2mzN11vunSBmTjSTQoxcRKOrrJQbhj+M8RkfmrrI7kUlGKBl5qV6T6Earv19BMtVO8Ad
/4ux3b5N3UWLynG7zRcuiZNVfrvDthsQYUgZj3G9HbjAfo1M+iXDSMQojYJ7DBwB228BdNKh76Vw
H2wnIYwy1PTq2KxDGJ0GXT+O+sisAwGS2VS30xb0bL/FAcm+uMj5jZ9VmdrWdo+/y1Hc8kHCbecO
H3JQysXNdheDyt9s06H0dXNoJkBJKkUsNwkYNjD3upq7av+x+16jCnG3wS4F8OirQ1eDaCGBW8mp
T+ogu0DDhx3+wCVVWB990pvcTVnl2NaBWh5ytl7wfrHvT94MM7o+E481Z1NzylPYJJB7kWeY1TQT
d6g6j7vfGcroeqr0XTVYWQXGB9xgRRKky4cydc8FWGCtnXw8nXAeAm/3eYsIS68O/ZVBx2sLDZBB
wy1AUeLjROYZCLB8McrohGog3VLg93/Z5tmllgwbp6YWntuKgjiQgWhrkgsEgM6mPDtzzgmKHhcd
clM06LDRL8g0qimAptz7PZtB5GB4vL/zb7fwkelDYl4sDyD2JAkCmLwyFCIXhVEDM93J/jRzPW3F
BhG0F/26HUdICvJ7t2AwxD/gQS6PyI8o17duV5w2ne5IKJOrxngn6tjTJdIJU7UM//d7qNkSiz0T
exY3y4G2SsPVlZ6espMgOgdpRFvaXzF+s/g5ykgjvAO3YlJzVKYqQ7wQGEh1CGtMe18jp6xB/JKQ
OEj6dQ8iZiZjmhMLyRiTtV+FdcVt0W0/9YgQ7+C8sMJOytlKsypsSMdZR65AZQzBUD0XSNnF/4Gc
bNTTjzzOo0ELhecOtlaI/uAl9M+bBx8pDXR625/cHyAXjjkk6OcdTOaRWmWhlIbNFk998973pnhc
c8pMUgvF5+Uht4p5L6jBfiOWR0dxzE92lWCRXDXyJipkVVjcPLQBIH4aKP869CtKS9Z8EBp3YnvF
SxCZU7bNOqSI6ykjYjpru+0CcRkGnTi9FKDonHo2c71E6dpSz5elHSv/6klsGwhZK26VUPimNS4K
ckpFr2FZh2gx6VrBEjY4K1X8r2H66x6d7Vs5rwd+Ms82+4nD6YDTck+VPMQ0VhSWfy5MatF+oX7V
uq4JaWWJae+RjEIobzdaZ3FYwBrb/khFZlnfv2gknSHYdHKcLvvYQQ+6friCLnwyhg2+/+KkNuJO
ErsQwg0K3bQcHPrd6WSteq3KmFQZnLVni2e+WwLN8zAeU7TPy0C+XleyaJ/jUbAlZl6NPPqZpvKm
AM5JX3+kNr+kUvRoNIXwwEV8uqohHB9Ar0UFFr3ED5dHeg+dfPSQX3A3E2VsGCcj8DEm+IYHGjtJ
If9RHWH5jZvUOQrZI9an7xd96RxTW8gtTCmBUj9f5fZDNJ9ohiZPzQvzccAl5Jc3nuiI4OSGSFN0
eYu50Xh8Nk/bngQWPOHsgm3e8PNHtEOJ+NL7JA0UYmIRPHa772fRdr3NTAo9KyC5tTJFns2fv7mK
s7UEIVsrZpM5ybYicQCzETELGIaTvYgc26pFF4p1jeNqrdBHe0IRbFGzm/lOOIPWdreUT7mvCluU
WbOW4YJe4JEQtoy3w4X6hP4A+lGtr8l5BG97T4mT/dQnyddZxwpUS84Lef5eiPq6NqIV5tVNDlcU
NXV8t+6AOmbpIwlhiosMG7YyGHOYTGKGPzwOM2tDA23MCJuzUU8NoC35TF7KyHSJXttEOvPlazSK
gmVyegpkv6L8R29JoMNaXNwKX95r/xt7yhy87/ieaOHNnrLOuSbU/7lczAyX14yJ258/AbhPHrXh
eJx24lEJO1w6M/wEDId4EgJTAxdkyd4swXJnzhK95GSMuS2V1KwU/Jgbnt30924E8i/yCu+pw7f2
u7IH0Bwx35LphhfFfxc2NeFn58paeNbQxYvrl7N+Sl3iWj0Rus3JAYD5YiEqOFX2CBy5CIF4w5Fs
zps2Vfh0jb4O8ghIWWx5Xe46jsTrSSbDR/ZvI2CoMBmG+gMYdpA2n3e4XaZcjiiPKhde5ER7L6Bm
cWbgKjdL0gWl13AfiHniTagaif6x+rLZVGCYhMBYSPNF0Om7Mp2N7GV56Mp+Fmg/uqQm5BIul3P2
xLaIMQe//apufGKG4vp+nD/WtBqfQC+HyjmqgJLsTMIqesADcXbIy2nL1EhgeImOlYw1D0va3oIZ
WPj4ZbT41nsCQh0009ix2+Yc32AcJqRzy5/cRNPeNCEMjG93asvKBW//B/HuN66uMTBbs785RQGK
nIWEcjqR2J9fZmPC1QYhleK7tIceWd+5R1BMGiGNZ/vdctxc8SjYCEiKDamoK882eMZDSMJGlxcb
md0/+qzi+qzR1OP+kVeQ2rrvzgiBk7b49J/igmC98DISPGTyXQ+eUqmAN+c+aVARwKn52U2sG2La
RM/nj4hp2yH7zpzYLqs26JzfoaaRSvwb1B2/y64KHIGhyjAbQmu7Zirw9FZE8hmPxcRO+NPXHl+d
Sjwj3seoB8hKaww20dxKXIwVBQqUxiZEwYSvfLZ1i1RgL0n2oY1Q9xrC1BJcPRYYJ333RoBme/2C
Kg7XoHWdZgnD38NvitD1/pEkbSTnjt4R9RdNvIIge1h16EXJKF3hvyYi+Yf1muW6gMYn+CTCNfQy
AxNWFKoPWKuIAViEKzp2iPVhzdILqvNscKZ4/65Fv+dYnG8Bg67c00t3vWYjbCH5f0GdrM4aIFHT
k0Q+48wGx/rU16qAln9S0lRrm3ArpMcPq21ZVx3bRC/qe4cBW1sVM99Hkt8ckqxOJiRFxlpu44P8
ecNV70Nz/VBmg5HUUV3JChaymfgu73dqstFGOewe9K8KrFlyYV65ypAhCQZnWGNrsO2byTwUJse4
iqzS30N6Me4KJuodS6mL24zt7FwP3ATTATF+0gLIlO9BvYZuI/CtZM0I/zV07EfAP1vZdEaYZldt
9XOSQXUNJQXyrNOW/aY09q6vx8OaNrTpLPToOreWQZsKdXaFuYvvkFrMkgvo9WvBZOOXy8KSFcA1
OA4zrDbHdxXKVvBegDd7xGdxFL64DX/nu6IrvSpXQJj4AFRKz267uUaZrDBvM/iK/a6HrFWpTcwt
7dIJmG0KWydzL3APl+PHpgX4idwOjtYhTiTHk/FSv4LBf5FCdcOoaaNutzgtslP2gSlFxRWcDcD1
Dy38dGRvRWnJkHVz4Ryn5kCBsJ+JUyJgI6+jpRrRTfTXnG+lxQMAe+nbXtxaPWOcamE5T/WC40xo
HEQ+EWKwj/NkkWbb8XOA11pI8oWBI38QaSVZH1clFfC3Urlxl7Ku0ytoJTb1dIu5nuygV7WLBFvx
A0qaRJnFTXTHj6zf8OLj2uV6RBA3JW0g8/RAZErW9aRcsd9XTobasvzxDY0iqzS/44yyOmOjhvjT
xrc5Gz0bE7NPtZa4UTHs03KjQuH9KtLHr0M7Nj4OCvyeRL+/AjkDKA3Ls7E2cvZuiI6DbxAqVBjm
g2e8t/1caZuM5GaUxje40Hd/hnlEfCbQpyON6CHnzzxuniT54CE3IDZ6l6gqb7xylHurjOK/1FNP
41JMd6wM5QcD5U1doGlImVgdWaUCIR4KXGJC2QXNTs7MS68y88yCSDq2i6aXM57me3K8tH2kM8n4
2mrUBbSwjOIsXfjg+CcCU+InA+2apZSOfn81y8pvICsSqgnf4DalKIVsuLoxHCjtaUsnYpTffPjT
pXIyRvT7fX6Xsn8eeuPF+k/v9+HfvU1BpnlNstAWDqkEhcgV+5kKhFj41/d/aG89Qi81E1GDYH8E
58LwYHUUXpVrKJHwlDCKgdum8qNV/fFmwMm0FXPF8mWGUp0MEV/zQzGwSxuZpK+LdHo4FLHkBQ2v
zefqQxSN98dSyhzljAXJ7zxOdxe5ySU/1UfwO2WC2jxscp8OI5+eidLGXhdzAr2YEvLuusoH+pYZ
Iop8WwpG1epPkx6bvri3HIev0QiXUmjNQI9ytpufHXV03/uyLJara/+Dd1dR7s++IAPoi5vD/qox
xUVLjB3iwuSPLhSN63b5if27RlR72JA1aIxJIuOzJouflLXoepp8/cb77xBERORtWn19T2x7v1IK
hP/BRS85VJjl1TLg5YOSmvwuf98oH1lWmRF45sutwXFpMf5jvCpokerYMLqoal5VAuZ+VDBrCQk2
/V8sIyj87CaGWBp/awTrpgL+0ho/dGdinQXsjvODJYPD6C0wvLqxJjdD/9MtgdPLGxa5ug09MjBC
tZvOOmZE5I7fvO8fxK41Qu7F82AkJbUGl2dJ9r9uVsqHX63+81qQ8qW+4lhLSAyaqNwk07YXEseZ
I4QcJm2QJfin15bkDzH/LTii6giOPsNTqD+lHNtJISUldYk4T7Rn+sD6nQztQh0mi6VlH+kZzSVN
8yh71tPq/MGNqvyVPeqeaYrs/5GqcUHyUjQwCydkbElgZF5yiaVR9jCVb7ro6ijkc2GoNstWHJ/F
gL1ORO/o/d6Gz9SyCDVXX/5ORo3lDcX0RZmu+nEDz8nQIGHIKfKQecPi9ZMsOErvM6lojeLzx3lG
7SQHgWaPEPRGjFe6lo3WT1a8qLJFrOejfBlWXiEJRmiAhe+VEazwr0aHYgM7g+kzgsq8if8k1vdY
hOgCP6wJ54XWArYi4EDYl8zg22Zayw0sEBJ8IffxuMwWJejLNfy3kIP4xlccaWWVUEDJ/0RdvFRw
PXlB1r3KqypVqLVHjvFX21r82SyDUonZGzrP40+e4nqgz2eFNa7ZrMLFR+AlUq4W2GD3s2HepjYF
XlASIaTTuUj1HxGN1MEkk4EH6VLMLLGxfc/FYxp8kI8cICca/4Vfb0aGTo7+UrTBqC/t+PKvLBcF
ocEYmQ3xPW2g+j3FkjRZKG4gHariGoCBUPUnq1qccejkYcBZ8v4L1DmQS8pNwpPgEPrQgebIhYtW
zTeCvGwjsX8u8Kx8lm9VphViwdM5cDv4hoWOe3mq7RCICHh9GbsbYTCml0vvzXGwtNt/95XG9/ZN
GqoVuBXIKDYmrAGcnaPHeKBPtqZeWt09a9giuM3oBoglxBhzFq1ot/IWju05Ykw0cvMGN3Te4nx8
bw++GQ70c25ffnu8flrcmc0+/zopfUFuLSl9S3jVoB4n+vZiLaykFG3snp0j2SWitSDVlj6ox5Fn
GfVx5Bq/1xP4GX8lwrdXyhhu6tvtHfLTqJfrT0RZxMGORGPnky39TXSng7oldFXxMajOQbMUOQUp
hfCaYXtFHW05z8vL9ujtbIhLd5dfce8JnWMrByaXu3UTGyPec4U1a/Kl3CqsQ5YGpeJNTn74pFyT
q5kZZ7eEi6XW69gvHL2lxBgAdOByj+KKDmVjfIoYRalrpJPI7l4tpiTqhunhKK20gecfkYPkHN7q
VN5Xd5uFL3tVCoTsIo/iMee85jlsWQAlHlfOa5fY03frzQ4Zh6jZrbT72HOqT2jJdOwxRSQsXx48
VlrcJY7hTwHF2ous3Anevm5ClgobqwB6/9suTkYxAfGOjyFhTBy+Q/ERMVase881d68+5Em0f6aJ
25rVkOwZg6Yzeo6tLvRozFCeJyC3PEvYVUXjfCdPq5DiDdcpr46SuUDTAapBJrgWcrUIIGECJCpg
3cWBK3Z6HJRR9Rk04nHaB5OQpZ5Uz2nGS4tvs9UaEoj+QRGyoIJpWMHH+48aAbkLk64uZ82GjxIl
SW33oT3H5S0+E0C3uvVv8Usj299eV6hTTN/Nfe9aC6vJuW5bQEnAa9SgkQjTdthN0gXehEsHdFg3
nUKzwPrOOFMAdFc0ACzcn+VzCqmTj3ldP4e0TADDymbcT5AbMm0oWfG2Eg+q90OA8ug0CPFqwSCK
ESvN5eayFrfZ3/LXyh1UZljicVNbjOGs2XUdaQY1hzChsGvml6c5momLtQ7gb3TXz2lDIFHl6dT/
KtKi4E0MsxCyHi+gazgS1eheq6SCAlwMQpDzpPzJyUmU/RmpeswsCJEwOWVVugEgFGNe1BktV71N
jDNSw4CdA6zH67YSnev6+xqSuZUI3xqVlRCSLLYo06Zy52xyFGHz0pAa5pzfD8h55Z2kK39B7pFp
ANCN3S6UO0+iJTvVr0ndOMufXU5Gq46XcLCWFCatKyjLzb9XyuZJAfgDA324ho9/rS+vJKSYIeCh
nc8HzAmN6pwa/a4aJwhKnohB2dDtTGmGPJN28bVWADeDfR3AIQUlldjhcbKQmazXp74y9OIf8ehF
NZ2o0Jaeg8ByXfiGs5q6J5MiaMmGG7heRFvgLXE/zngLVmjELo8g7zFsD/J2L6e+yoGehEEUZq3z
YpiKkQj7gQ4hZBZ+rSqyNcQWUkRc/iC6Hvp7qWRMZzf8ak1GRMb1p9HTSJEWe5Z2PEwGBujmNGWX
2aPFfvMFEs/OpA8mWe9MW9TTnpTBmT339Cc6p197RH45+NuHMBgHG2Dj1BRvKWld07ske0rghMHt
+Tf4063lHb1pBkX0Sw/C8NKNJU/7ZTf6zbCeHobUsAoz3yTKwe/0cMcAXCal50mAvmiSNKGcGPgt
XzIt3W9Bq7qEDePS0iYW+DsrdcjqVNI/McTH15TRRXj/V89wl513nvKOvUoBFN9ppW6NqMlkD3qm
kKTFybnAweUrbTN0RsoHGmbXKMVvQcCx9EvDjA6K4JzGFy5b3ogx0Zguv6u8rIypPnEtHby4t/Qh
EslTUG1GMwHDrHidXIngAethLtZFkRwntepc4D8QMaF9oudemi2VA43gpJn2VwbL2I+gui7oENDX
vJ6e+1m6Vu//HsJPUGtAnnWRkMtyi5k2iL7LIiBUmmlsbei4gu7t6j7UZ1F93Yn71mEdhVwy6u6D
mxb2JScxlwqmYSYVM4oSnhbgzIA+U0XqxgblPyRB8l9qR13snvX0jXflLEsrG0UM0zdLtJ5oGSIx
U+pshbYsR2WxB73fvMQBsY2CCpVLomT/bWsNzESqUjBKc3l8xXQ6uJMuC4b3NT2qzzdHWXzDW5bY
11Z7stNhkNr5f+Vua7QjQFdxzBOFz0O5EO9tr3SCDuGIqKM09y9b/c6Y7jjKj6lwSDTjpFMU9G+9
nsBL9eGXZXcgtGrfve1/yJjsTZz+1/h7rdo0LoeYS6cTpktWk70QkEOPz2XB1R1Rt+L/NThx9g2t
0uJPiYTKrcGtG4UeWx6SQG4B0vqlkM4WtCaZElY+4SRFiUWcyLntMb5P97K2KCEUWXAqvR0JYHm6
fNnafEUWRyzULe5WBTZti8zCUO8eL5Zq6bKPC3e2mW0pE6xxP7HcQ26cYsLTzgNCuBPjZBa14crZ
m/vnrKB7U0p/Y8oGzXrhjGY/Zbsaf2JwYbkfJEBqGDIPlqabaxsN+671svnkqIkd1C0lEypIIFm4
09P+hHT1TO9GKs2SmAoxBuZ2o33BJ6oyl7PrT0JEJVbURTc4XAugwj2mMbWb75iqZJoXS5BiDhLE
vvcWsdV9uuPItyeARvgVySfTSlFGn55lhop44gUYO8UM4qtA1+an6UC0jE1hfMQQZ+r6razSc0K4
I3l6IVBdNkKV238OMp4B/YgJhZ86t2WpPOa9u6BctKocik/bljHiMSSAsJ70yzvY1i5qhH5mXlsD
wn8WE6T9T3lbHK9DseWgiEHj5xQHNcaNdtTlCeGk0qyDJe55MSDaxhJnnxbHgTOlQS8Vupi0nR3c
XAo6z0iElxkVOJ8anM+YmAEQSN0YH0d6QNj048iRI8mWjKfdZM8FRBJ7fxy396+15d4pPTahGA3u
vPY3eUUGGnBFg/8y+4P3OVEUwE9o2XQxt/3R0lRgZjD1QaZ9izzV+rNucD9qyM26DCG/uUvJcBo3
YQUIxOCOGIhTFiEtRL0iED4/45jpNHgsI0dpe2qVjyfY93HxF97lclXdAM1q7Bke3CkHQcv8zQZA
WwUMO8f7jGp9YUfS6dlgucCl4ZKFdr4St4tggzEwW4Ve/0NP5FN+bw+coxeYE0A01NPJNfi7KKeS
B9Ab29mFt7lbp1TTlWDRXWR4jW/cn0tJ0oFujlzV2jhAJ3wNCy38bazQqvlJw9CHFZ9Wmuifstmf
IkY/zvEOMaSIMJdDMx905Quv85ERfOpECFmUiD3HPaobfTn0S1jw7HLoqvifKrAPcmHjRzh1eMbN
2WfzoYWo5rnmxUYG5qMjZDJW3hIAS8OD+i18zWlLdcniKINGHA39v6AFpj3/TRiTVyGjr4mBqqjt
gUyMMcWZxKqvcph3wDxHXdRVaGhygsJqcHQftXT+RRkhPx3TUAjvHg6Fp6AksgJo/aBvYosVjvAV
MPn2WPQkdk3LnXkNEHrdC6G3ol7KUFhiDjtYAtWfyKM65wgysZbWa5EblkFuqkpeRYC9+SgRCbii
c0io01srp8U5q1DlbOx/e+Ag1greNW46z2ENRVUkFG6NGNezP5eCm1y9ZXnm5xfSUxcUD8A/GJhe
sb95LimaT2ny5UDuPrYw4P7/ARK2z0OY9L7w+GmaKJH+j2mriyOKT1psKx5l18oHncQUJ4QFQbSB
ZnBzUGaFUOsF5HWgAAlE1E9Qd96C7R1DVyFrvq+fyiy0uAq3dpsfNi2iZB6mqyX3OnhErxllg5KQ
ZwDpX+DJhZG+uKDqD3uEVG2Y8Z0KeM5/rWdua9bWO8V5hS6BXU2Mlggf2jvbrkTqB0sRDqTv59J/
JCiunb/K0rGcKqsgkEPuFk3/gbh6b/8DmBujRWtOlrma03K9/ZIF31HKRY+o+pYsC9hsXfAityVF
+uNwA9qQ3ttabTyUat295yspQNbHffk1xxB7YQDaei0ZnIuyKOvdrTEexureVicprMpTDl2GCSSc
M3TSvavfUKFzPyNjiDe6ARUan0dmAWjJSyeRNb5FIwfVG0kBH2R95AjUSbVQYrHIPd7lMIRIJPox
yDV2ASfHMD3rLd4EIjBnIKAkcNip/8rzkNicVk3iR3KmXUoIlM2G7HD9mlCP+ikpfO9OY7td0oil
pLRaS+GIib/sN4iWjJBVl6Rd9LHoZerXgGyF0vk7r7x7cSYLksnRTrGN7APGwcLbCYETVf3pNIG1
vjOxVzWBr8VgV5PF2Pm1luiad5Q2gxcu/LEASTtzHXyufWhsP50MYCb68mpXHkWbiaha7n+yjZWx
AUW7odRtD+JKxVGNvJQ8ndHS+LjpR/zr3BEIfJqDJqU93YLbDtbqFsd7ZC9tKKvavEDuqSyxf8Uj
uBwlf/6ii7yLN0zCph2PihpyFzW4k7G7PnSGTX4P/n94M1C9Lovmuw4QC6uQMqLv8YMNeBlDHD9u
y6P7705sRceKvfeEq0ZoDpR0Q7DA1YEAbZqX/fu2FKMGUyX3lJKwljlNAB8S++pSMq1EMZ4jOCos
Es9RXeI2ao/D/n6wW4dWcQPXa53GqrBcKgdYdZi6E2OysRfK9PT6XDJdM54FG9k7uU4SEhpKdGYu
KKUUnYkTyuN74IDcXeemCE+QfrTalgYEE7RZetlJsm5E7hCSr+AkFoxS3NYDCuM96CnDykfuXpkC
fmANHGprjWEI4AmnBnQitQL/aC79wOukCrKLABw/QBB4U5lTkt2xOQ+hqFa9+XrJiktJQZKrfGkO
FzIbS1b3A8v3JU5+sfek7fZkOR5jo/+sXvi5HEV0uaOTc2YseTwUuMPVC3r3LXLhkegBVqDMy038
wNz1iPR8H5KedgIm7H9CbUMvTeiR5+XNDqGZHOgySHcEEcvCECaOHTJ17a+I6x88ohHSbzc4T/aB
4eEN842M+8jpldEOMuvSV8F+sNsmdZHvZMlyixd6P3atpn9vnUsA3VGAcvX/aAFBLqbLpL7RrtTm
oL1AD5mpL2U9Buiczz0b4VDy4BAeH2gMD5+uotnDtS91DBgPPZ2QvdzZ3n8aFVNawLYwMANPsjAu
i0RFBTtKjdsM9BJmBNGsfw1fO/JXZqv3ozSR6Qj5fm0nVbBMxhF5V7NYeiq3vOMxHBPsfXc2a/oB
FAefw3wTqrmfruMCjxtYKXv5i9ro8hcmli9BVzzfS15nESwimlepLH5LK5yb5RASR24IJSsGBUFq
hQ//RX27NQHlEm1EVRpp9uSaCMSTxCrQls2FnSAJi5UuMoovieND6OeiGQHeeMqWnnPEYsA2SAIU
CHN84Rjjd/Zq62xDK0itPo8dx/7JQk7k+IFJu3YzQGmAzJc8hYfphrPHMTMQCd3kdR7BPxgr91uJ
PXy6vfMlwiLad89k/TsCjSqpZZ//W6sU+nMoxDuCrRUOzWS5NsQooVHuOZIq2YhjLKlvrGb1KPXM
Q6uGvPUwUvCwe6TGc1sdlBa+gTJRDIJgFexIEW5ceSGStmAzTFzMArB0TRjJOqoo4Y6RJUPvymI8
5WThMSeOAexu0ugOIKHaJAOowSqmls9daICDEEIvpxoCbX3z92LOb9sMvzSTrVB+WZk0t2x58A5I
mQEDToGmA4qZIco5QVI/761TJsCAmEjNvcFspeEYGunKa9ac/uR+xtWiLieweSX9/Xd9SvzsoE0o
GE6qiXomR/C/g2pGhoZS81+nVh5kupnUE09JyRkyMQ3fYjYCryxtb8yfM5Gz4AQ8vHo6n+EnR1Zc
FbCpKmf4Zs/1ZZb0h9SE/KQ+qiRNefuWHUYL0DmGJxe7zaVjnQV1p3FcB7X2SLEAdEra6/T/x2vr
2BRbMJgg3z2bFwNZ/AZKxF+WsHNmag46tvwvjSCKpEF+cmM5kOcsx6q16yhXiTwsxlKbYJ/ZpNUP
7xeATHc/vUSG0EqZzfRofnb9kGp7ZiMsQ6Xl3Vmn7ZbLRvFXeGcbKZBw3nRZHG9yAKY4YFZ6luvV
bmdUvl/kbx8TOLYD7MDjgnjfGLSneTrssYwQcSAkFD/E0S2pJ820sqUvVvu2Rz3ptTtqrQkq44lG
6N46DnRvJFvUUwsOaRQGEEIZAbOfJ1R8QNfXkMLofhQlU3ztZtThRY3hiukC/xs0Y7/gYraA07dM
FnTRP7vFn8T5JSZwqHbZlETfOsAY8okt7l2e4uvwrTQFOpCSc54KZ3AMpQ+0JjPjQRJhh1WNMcky
lNjWDb5BqTSyrmTf13nfaF43kFd0Ooxti0mkvj21vKKMARlqjUtYZK8uHlA98bDAV0MDknjkfn3+
eu+T1UEMIXBMBbh+9dequbpwIoxmJpqDfKqv8r3XNLgb26YCNThvng/wXPOmSvrqQAlIpixof54O
l6SE+gUPyLUIb344zrpYztoPvYx0ZMXaucHAnMMAusgX2Y5KDwili7r7j2g8go1HB4e3Go0rZzit
wKRBAiWdqNDoSN2VtXnoXQhE4HyS/cXZOKT79Pf/icLOE5U1ff2p2o8a5V5RnRmtJzFIN/wHrU4E
bqZDM/6pBR3y5dnRbYCyEm/KYZ/HC1JPwPf/12rUbBpDSFfVNGj+PH1iiU1XdQrEqNdCWNS3qv3e
CFq8zH3I0FeLWx09omeFmb2o6aO/gGRtTpSgvX8KKp/M+0y0iyCvxoJcRRlGlKP6desQ1Qqgl7R3
4b2bwotfxC7zZ9h3TceX/0x6DOIR545Z0Uh2qyYjt/7mjS0Jm/e+F2BQxfEI/r1PYoA4FfDTABbD
jMWoGq20QIxyDTZ2SyC3CQVcGfx2qAbzmeQlCTE4JF+BeS3QE7u2rxId+VzS+bLe09qXSZYx4Aop
XpMtEv2lw9wbNHZq32Aw0U8S6Ok6qq+fKjkeh0G1EdXZIMdGr6XID/K6TUTG0NIpQkpfLLiR/2Jz
JAVuLlItMW8reD1gqYJoMwlS1k/qrqBdHwL7rgH3zvIzgReT0VJ9nIgE3yctlU0a6HmquBksPeBT
Uas/QUjdWTOUc0+vHRkE/xClbDnq6f56083+MibJNtnd0tBhRPHdL8cC0vhleq3bfIKHaMmlcySF
a07o5mn/KJoZ0ziRbxHSdElbztfVlKICcRjH3JkoVaoccHAi9AmtwUCjhZqtPj88z/VKpucUk5Hb
8nF5hNi8ZPMTQFu+/F3qS/SOF4pYN5k2YeNhDv0e8DYjtqf2Q8wTiJbb2hUKXQpPEf2aFj66D6Ag
1Sb2xagLBve8xCnEYBHYf1aAvkjz+dzs2hijSzm/qfFQ+ZPF6PnIs/dPPQL0FxX1jxSoJsdyWKTq
R+kib0zn6naKUlVu2B8ZGaK/5b5VJoUOFaN4jvsZJ5o2BquP7aAmf7eajT0mmLJv+FKGIZc6YKSb
OKjohKly9m49mckEzFLyr1F19wx2FVN+qZL8/mDTITIDGNvMy6XYxm9BqWmZdMtOC0QapnPCAuBH
iWG/q3qrvcizLjLbNHic5xfPi9bMuC3HiqXNfaV0XRR/lllzRTNHBIQEwFKE+xHzhCZh7XENNZWC
1i/Q6jFsws0rfoAWPJ2dW0GyDLR8BFDR7jyyZ7ugEsZ+FHqIyRi3kYOimi9D7JhZzicpq4Aju6QJ
3wmejTudUAxfPnDGshz90BDZsu95O513TiLERAs4HlkiwiRJ5Y/hyvJpqPmUx4XlNInAE00hiZcP
H/AiISntmj+GPsEV5A83paGXZcySXeB+dtwnqQ0umX7N/hBmPHJpC11ZpikPkUZln4SEdtQEIlh8
qsjtVUkojFsw5O43DxWTPQ3fiSPI820u9N/p4bWoqEctmo6yVp+Gg5eEnZf0EdAy8l6XmxDhpjlJ
91mlK792A/8cbigpiaU3hTReZZa6N1lEGmBmVoqoDwfntkLiF1ccSgt5TRH9HFNG2R1t0EV2jS9r
FcJvAKWhEJKlB+ySULAPs4FhI7Crw6VWYcroD7zCIMGhV2bGWcKGj8lsR0Y8ax9bOXsni2UGIvOx
kUtVLGNT7mdeQ1g2OGujOTv3NOOsyho2GXec0EL5B2YwyhhKB+80rFytsyhHvs5MSdCfppPXLuko
gxxxhzNzlEzD77tdssBbfSrvTpIFAnCt/mVj0hJ4eTYv2gIf1YqwkJ7B3RSiklmVliYWBV93vEw1
gFlDUxEX+J15WpK+TB9thAelA4Wbw7Yo2AApTPMNFopsjWnypIky5yxnfWSlq5sYJ0Fzxrzm3U3R
2ewF+3auSQ4PY7+7k+n+LZ1VYxNPDAT+L37xgfg3Kuj/o5ZnQcZ3l6Pua4DAXuZXImjh/Z3deCmp
q4PC3P/Jch9J+/MEp8KlLjtXgItoh23xOqWBG0OMpDpcFVed/YWH/JtgsOKPkvQ6phrcXvMwUoj3
PBvkPHIV7X3DoU6s3E6g/TgRIRJ+dx3+6DvxFeACxR60+YukWIHBvs+0Zq0MDN73z1SQIIGF5Z8m
sjFO288VkfkYPNUg06simDOePNGEt3NX1zsPwVW8nlhb7y+FL17HoGpl7DziaUu0Yn7O015SOcmH
mHU/c/phJujHR2Ty5XkUKZLTmxevypivBcwQgdbyGVvqT2/NRQMNSl91vqEMxF2Oj3Vryf8yf1pq
WID9v16cyxTmyirTw+Hz8R+f4bBA7BwVXu6WKJCcrENV84mYYvzQ0/VHWF73iUTLCutmx4vPXyXw
nv6h+cntHm+pwQUD6sioE92beshXPnPpa12YksPOjWZ9F2WzAxl8Jg2FAsMnXW/Dl/ZpBYhkL/SC
fos21iiAjG9h+tyduIwkkql2BIv3F06mHUbOq1BGrhzM9gQ4EzzHFCgG77kDmSEsjAw1nBT2eqwg
T9hFSDhWWHCK1S4n40VEhPcw9I53b69nveZtF8/SFbIwOmk0Nr0XRzOx/bwSKZt+3hR+5o3Y84Sj
z+pYRdM8f7K5q8IDtzE0UBKVZC8WNXC0cJxBi0pWv628JW3REec0y9kMmxbubJYbaJ1/nNZw/r0g
NVjNDb2+8xkJRwgLVaGyahAercKgDfD+YD0e/QEg1BtvzR9aEpqc6Yf1cV8EmwL9EdnUdxcJwFxF
u8IOAE0mANX99jkHMQm2oKo4h5DBY7ae8Ep5Igg4yS3nMlYkp3AfnzYm6AwxkFWWiRrXH15ybbtz
ttOs3WE96cEEeVFr68Zagpy0f2WxyOtVeuDAwojaTjOm3VNilZsKTVXYEPsRSUrwsHAix1uOTrrt
qG7yJvS1tnolt0erAiemvfIyeRkvONP2o+IWfvve47Ost7p8Lej8NooCO2eCU27IkYf8EtegZNVQ
HoyLPwJWi+DK43dQUgib1asvzm1l8NiNdf4jAkLjzjSkEq26VmO6fNLfBDdz1XQpjXVQlcG+yml3
gbe5kwe1P09XTiBGkZwzy10eVfBqiIM91AVHG5B8K7RatP4Bbr/YPkF1xm59osjWnISwY+zgC/X2
Lg6dK4ygdIFEWPvnCPNz4asmMOSbfhWwTOsiLB9xRTDZoRka/lte1TaxLwO1PABrmRNWULv8zrob
ATIRksNFQ9Qo91t1OXO1qHBE6MDzI2xlRTaF/1yUc4A902dvwS3ga/457f00XYA8mnLq38QA24CF
U+tFDp4VAyKFYNVYJ54sxmmYbYYHK11a7x0dYD2YV2JB1/o0YtyLKR6fa1/xl9ZUs0XNWujHCPib
/PGSfdBJ0s5NlVtZkK7EFy9D19XdqGFPmUI8BFV8/rSa2i3LgMqjGRwCxcS7cztFZqe0WvdEhxhc
W+/3jTvsrl/spHRY5A2/5JDlgeCoR5j1tBhTxI4SUA0TbSgQT806QrkJxc3HJgMToNAG0LAkSyin
SXfQBm6WeEYEcnV8HkbiExalgqN0Ke1jQziF1ezvXtCGFroFROZGi6e3quUWyTgRemHbKqGySV/F
0RAHi1msWU6OjDdUlhkM4t35Lo2zo1BSMbRH0eeinx5Q7BRKm7B8LlVwKssdX3bCNL19NPGu+X4S
lmWBsPPDY0NiQw1SrbChVLzzT6kN7hZiUSWS7RP1a7OyYUybV3q/kCOnxTwSmlnJwjRPrYvBbSLf
TTgX6wHDatYC8+mrnFSPtl48lg1aEr+rI0mGp/GXtIUqXvn/axlLN9O+oc/Cq3E1qIILjE50PmPR
yeSy67ae+wW9eUbWvqMT+1vRXDg+JCmwwcYy0QksmadayC3ystqGJiWi2yKclsfVAFf/P8S6Z5z8
lBuRCG7nxYPj7sNlgbkmVpyC5fXsxBgV3FfJIyDu3mR0sB8vT6Nf47y6Tfcn3T6OyCqI0GT8cbjX
AKPDddZyvkAj+eHnW2wQuGG9dbia97ecUHrlXU4iSIWMbBR4C8klU7pWGClLT9aWo8HmamTSKXI7
OOnJTUquj2hTHcGjPxAt7s2NCAf/Bx75S/ORRIg16T5A864xaS7B5x5LBIsXR75I+o7iV7hIr56z
uhrOy5SETkt7Pk/645E/nrEc3IOLXcr1ssLxbTZRRTDTWXJnqk8j4dKJS8Q107/hticR4PHLtK2Z
lw8uQdD4IvLr3NXPr2AhD4fzFLa1BuZhcD5Ah5szqwjdY0ZPbG6MeKRJJ9S8KXrbVttlScILWZc8
4KllD6GuGhIRYN1CIZGDy9LNdzxlzfFqfCLtjs8bdxH6uDiYxkg1f0SsiMgPuOcssBGTGp3dKAWZ
Q3ofefoaUD2KBgyQ1K1AespnxjAb4Zn1IUCL7OjRpv9925lx1WWT5DS7w3MpyPRIk4+ARdJGIjz7
ArzpHSWGtNayV3lEMYUuX/nx8Q8MrS2GCvkHoniuesGXM1j6TZC6KfVu8/Mxdso5vTp0mMXAkHzN
p6filayjOGShol3ee8jr+trDYuo/2HaMgXnIZTs5nqJ9zXbWTiTU1U9cmWe1PI947RPk0kDIYQSy
F7evWrDtrV9UwYvJAdUi3Wv5u6d4rMV7aK8+IQ6+9yv3ZKCxmvh32iVeyvsPPcGTunl8cuI6yecc
Io4LbQqJakQtfPcjMj7PxOTSI1ihYpreB4HrbX+KIErT6TrmTpUeRgz2K9RcgEErtgDKk5cIh4Zp
7ULivHe4yYmFHg6ofAU0oYmhcS7Y3C3r7KPuugd1TRXx+cyGBNmXLs8VUkT+FsWRLwtd//6gB2hc
tPXG5A1GN1irA5wzhfnsbV1kJ5N3wvZhi5Oj0PGqwe7LZvlI7H1d0jgu5ybWiiA4AdIL/b0deRq7
ioTp6UaCQQ7GKoE1aeMC7GF0X2Pnf7OzHcySm+HWLUSgTEtnfBVtcEiRxDc+naq1iQAV75w8DgrR
a2WjN5mvWcuk3+us74FmSIvlQL7JjswPIZ7d3PT/vLqW/obNNh2NclaStR44WNdRPLCNcEWOvbRR
RFo9foF6JkfQqKFjFMb8lWK5zn+trpF0ZPkWPpN+hVc1FL2zcDP4i3Nn53SzO+tsJLT5B8CFkyzJ
LZ0fk2KyvHTz9+HLhHGZh2d3gEHUe6Pa+9NTnOR3zcnb3S8WWUhsd+7ybgE2W3bwHZNY4YkwG0Vk
jHFunN2/bOupnqkKDWDsMu/r7sNDiyNJHUIhORhznIF7q6D6xHn/oKQ7OBTIF1hRnT8o1DbnQTWQ
Mue20SKIWZVI6Png2zvm2tyN3nPWRtGP06Avmkd7YxHQVz2EO4gIbgdo1d4WQOM9AB4ga+RYeq6K
2O/lYsTlWOCjC9kD0LVvfNHs6RttzRzymW1NcSJISeovN89b+a8BKPDtiqKsj5mJtCH52tB8QQvQ
9rl9sxE0HX4th10neRrac/96bLCbcBiqQLHS5dFq4xwmsoALXOvxhIlueerIvRJdxiXbULvhYDiX
7EnY3ITV8/Qh2zHk6M/bD4uZNXjuODtJemLVlXVl5qYIG0I/jBTg8liqtGFUDl1Px0/yU9L28Wk8
1W/g0CgkaJFnDmn5Oh/ZO22AhGF4sB793QDiGCmTWVGwLWG0ZHSi/GUBfticTaMjeyqGDIa9vzR/
fWpSe7Cm4Ew/9V1xfadGfu1uczdddFac8mFyL8K9i26PoWSkpnsuUrsOezp5qNSIz457frMLVTgR
lIUJtb87nYnawNT/xJCdKUbkTounbTVZDuIiwUVxFwZWlD5XG0mVpTgsekH1D7lwZOWhXoiUO33A
aUt0uokiODr8a5b1djI0NWAmGB2PQ/ymxZaZ/bav7/WC6j+I4xfdP8O756m6jymfX3tEbsaYl9hl
YZcgn7xGdHzqYQZlUWeQpfKu9+xx/vCj+c2cGkP+ws8DdAU/wAKx2PwSPbEriLEWGKdw6T0PkJKm
g43IedPpcEu+kqTzJ5xCYBiPRl8tOjw7FVZkk/WU7uQdEGoUNm09zzrOKNhd6/FH/SAY2lHnsTSu
V+jB9lSN3gs8LYoy4WDomKl240KGJ70d4qG5SrSvMYVKISIAUg91zZfAimrnqfhpPwUjJQv+3RTz
rLAVd5pvPkKGpS95bKPdJebUXWGy4mPTHOZZq6axCAE7t6JykMNGYRJqxFPyYsEWJrCfray0pniF
eKV4EuNMirvHlbj45k1TnmrDJmtvLtlfM9X1//uWLMLjDI4tRagdlflh1Kl4dXrLX2C57E0bAlHj
jl9JHylP1wcAJCuf7My6DAw/S1Zc8keCGaGhXMO2KvRuehmbUfAgHSDQWYQBsWwp4gBDk2BjLobw
MQMXD+eY16LuuV0V/SibhdzUHylEbXMWWouBnHFW/3gHC7KyaEvpY5fUsaBAvzQoULgF7bweapFj
HlWICzPSNXCOF7P6rKREd5b3dguxn7IEWISsZ63Ey/rcH29UuHaZlQZiFWr/3/6OpzgpMjDa2+01
x6q/QMBB/c446VkMZgCItFkXncxRtwNqSWLeuI5sJ7312+zmDcCMa6KDmLmUgHWfHAWi/BceeoQL
LKPb5Tko6cupJzmdz2LurdsUbrZA/PZVts8FZrPcQRIkEzMnRAmKnKJbvzH8rd4CQ144RIZXVYx9
vNgFFrKewiwVqUlAPza1lchVstcHncOd5ddVslrGRApQJcj8BTku6AS5CXdNOaufnMmFaLECwI/D
L3OEToVosMoVLRgfbQsYiCT3kdF5CkITPRsN/WVX2MaBGlbuKHosJIadZoiA6jzNXxaN4tUhnSoS
4LmyTyE+EkBBiJkLRude/ouOXOnmYeEhzj3XD/62Ue3Sc44bZYueZ3E0LNw7Vf95RSjYjzk78QCi
Eb5ZpRVyyHQYG+JgeS7Ak2tVfS3rF1IYGLD/gswx+1FglS3wtwqghwxkRLFF5Qx3FFhCzYj1+Cz/
gpWlWRJzpthYETK3HJf49+0hoBb+VzRXhVHQIDyjDe1RI1BBV93sPM13MPHKsDRTbtBne/k50A7/
HboqDw7eCi5jksj6UjJ0cDX4sFmgvMfm0nFX1Eo8Q7x1UWPo4mDieX8MoiFMtlhyQCRlZgDAVGcl
ncGKjTQr26BlkJOhejv0od/9J4AYte8wk/bmoeAKEMSsJV0ElTz4ttGqeKcv6Bm/QB0dhYczyWEt
lvZr+8L/TaXP2Fe/dYpcE90lWSi3+sS10oCCxtMCKSRT+jKeNUmJxazUMJLgetIWY/C8JOA0ayU5
iD3R9I6+eSPrjpEb/Bfqrgy+AQzGeGTcps4jHfufo0bfCQaGG37yfs0goCgKi7CHy+aSHDTATzfL
lun///B7xLtlTGJVdEtVQX+8mTPz3yYVQLU2cn4FdhM3KdIf1vyHNSp7cWck8x3V/hIBcoQ1Uz4J
nu8mw18WLD3GY9d6q6lvxy/P1SAKOfchP6e4/ID3FrsunQ6qdczMR0chbeHCN3+HR6/Xj3rlTEFo
qLHPmMQ0XyU6XW7PfIzxROnwdwtMzS+5TdWf+ax+ndndYnAhNA6JjCW5wvOK1fmBuJonVFJ8cO59
4UzJI8xhMyOVj6T51s7P0vkGX5X8hi5E0xuVAVpMe+sXT/keHLjQQD3JweMVXjkPNt1K+xpzabmX
SmxQE7s1a4GXz7bzj2KmPVH73da3BF6Anm6tSaekf9YbVPdbp6qCcKRR0vHFkD25UiNgnvkd5bfw
kEPdA+36dOc5iSHKWPIiplaNcp2JwJ/b6eM1TmM2aj7oGD556b9yDkOK49vlyt+y+lHGuBI8xvHY
miMbCZQWoJu63YZRtsJuaFDu0fXImDAsz2ifqaSpT1NWPuq4MA1SvMDIweBzmfKme0Ky5r1yYXNg
oLWWAYUleVu2BtpWVWcZQc3BGaH3nSb+Ol0lT+SOr4u5hAnwTFra1UGlTHLhQYnTeIXWNDHTVymF
7uaaEUEd0rtBcVaA76lW+oHHkoyqIwjS2gJXQaDyi+kwwtQPg/6dbs/1MnD8s0Ich22xvyx5Ln4j
5Fgo70pKOf1XQ/3HCGyjaNacaQIGbpZVYlFigMZCsqCckpJVkdkkngzYgpan5GK+EKeMhCNU62gn
+lfGleCiVhjPIE1w5sBxQ7efxg6BhltasX9l77Fror3pYANTPEPYg1v4DCiX0tcHEsZbdYQ0ySIz
sblt2/yDtefUB3G+7jI1PQB45yrBveRv+zihePdqtrkBI01qhyQe9pvgUt4NxIFwXLNbCteRmvrA
Zv90fb4LsFZ2AWh85rKdp0AWElRuPXqQS1u5lPxzzKa4NWZ9OD1uEnwdBatQZbMOZPQFmL58OeuE
yBOSl91/9Hxd92ouwsNeR+OvNiw6B/TYskKqeypOMjD/2sbVkTistadbPXzghZ+AmssHrqwyLQLn
JzBpQK8caMrUghpVUnpFFF6uxpxkGQF9ctlJMNOOa64nmfl+eSRsYL2TGUqDuEVjzjxMtFTqqf/2
ZkyQKtboO3jOyudur5F1vleppD+Autdzh9o4+8LiHAMrmwBBF8DphrLAsFmVMDQBsyyfa8lh2USl
OgjeeWnqmtcR/QvH6NoOoY+DLzVQbnKJIsnQKXmLVIWImQM3Aq/V5c/1UeB+kGAo2gWTUZY8NCfy
VOOmUcoWTwJZlgmszva0L4xHM90AcFu3fGMEVlKlp/hFUdWhK/+Vi4XXO55P2VCC7pXUqo7ySrad
9xyL8ccEoAXiSPtDRQ1jUT7+CjPoILbKZlMnATsahss40YeMqp/M8M0zIutLFmVKQInj1WsoAogB
rs/QZ8kpkTLIFS0MVJH877ptTVjv1Ths6Ldrk8cjl3EbA2pFY9s7yBH4f52P3n9lYHDSXYLesJEU
Yx6yF1weTp3fl0EMldgHjfPHzZ5BRdeIUVk4usMLBFUIsKyTLzLiGlzkaNdUfSCCmX21oL1HcJnR
L/CyvJ/ixeoNZW8hodcJgCsh+k7W+TBJJJs5g64PBq8uMWrSz6CO3ecEpbSH51stpVrFErtEA/Ti
Yg0S+A4L3HJ8ccaFRjPEsDypq/VAyibcbU92bAi7lF5ACxGMmy7oKAOQFdDmRShetqcqP87BeFEc
2yccHYz35W8IeJiQ9GzwV/jpeVmQaLFKIlXW5DJkebRlJWHKTlZkVxMJDTea7UyzRLrxVsxe44Q0
tXLQHgySbV8BAUDxXvKNi2nNhTNQRMjO8UfDBZ1BQ1xCK8D7vlG+wIMYpd0i5BcmCqsiVOHwDBPn
mtJfL0HnhdztEZzYiCT9BexzMX94Sgqi5sc+OP/colGnT75wfOCpXv+pNhO5R6ekwLdniFQ5crwg
yCQ8R+fLTCRLE1QyDb9dS6CU07npp2mxJxDJBnZZuGZWYH90EjT2luIFiiVPZp148/mtN/zXUawf
0KqaJ3MvfmR3bBsISjB/5kjrpP8jqLLU9dl6UlbMDv47xAwHZIgo9u2/KIWtL69cgvzAM+NbQoiO
qUM/mAdoKnSOk0hy3evaNwRhWxmdCW+pqXcRU/WfcO21SNHRF3VE4I8ROtJBlh35/sudawB7pMZd
XVyaNb747GqWAZe+qfAvvqvHzL7/s4U6A5gvvERQBuIkVoqIXwCX4u56r7FWamRi6909QViz32Q2
teNeHh7GWdyCiZr76G4YDmpvvuihZL90gc+gASwb7hSweMxt78mbW2U2YeNTk7WCFX8J2t2Iji+Q
xiWe//bEbKNo2Fgybz5nvOQLzTQI/vU3ci53LgGqxgBXkcfFuoBRsg8eFrJCmuL0Xb5Z72gP2jR/
T2pJGsD45wkOE8rKGspVHPjJ2N1yoYJOMHZIrdRzBq7F+oLkHEzFbSpBYchwJrpr+xx2swTVrVYI
Wu8qKDXeUAybd8FFd+0B5UGp3c3Chy3v2suJeO8GUMBg5sF4LL9Tk8ykPAF4FmYiHYTJKee2XcJT
uFrkeTqOH8Knx9//HXJNqwMyN8quU+ePp+WETlvnJl2fIZA1ksrGfOk303vEdMfMUiFgGk9RJwaJ
VN7Tyq9QIWZIMYCuDCR7yv9FMdg8vkU1JYMzWdLRtkeoZNuI10pf+fuO35kJOHIvAGaa6e31DN7T
IpcOkXPKqg/HTKOe8z0CAGGu1IzTjopfpXPQQJhEJGjkZaWGm5w0Kr9zJPFhE1KlJS41n2rNI7Wj
tzPt4Ma/PR0faD7kvcdU88B+MwZFrjIzKfi0Xsl2Q96uzM7Jg/ZRlGae7QYlGHfHO6pdn6lKczV3
iUBwwdu1irGZqyA4QmWPwri0v8GV0SqWqotM9UmvxmKtl9JsJaJoZZ281Fd1vznZungTW3bREPTg
SbZXawvqq/nNpKvE914Au2E/8/nRnp6HV8v/JJPI9NMqZlg/WY4yd+t4M8340FtkY/ynfz9XXcUL
UXfSPgsd0/IT8Lbyv/WQr5REY7G1GrCgUzijIPXTdWe1PpoKhlSpCDZ1OTYTd0b3a7mkNevnf64j
hqn4Lac83cL9Gieuzjys7ZHtzG/Q+RclKK8mglIySixO2qBZrwWFcZ/ZTnlooozjrGJ8IG5GXGCx
N1OnmsxN3wHx3yy1ZUI4xtc0oD6+qiRJ35k3pNsGVWfNefSizY0ka6rVw6iqIZZfjPRq2QMbFHrv
03T8nj7jIZzlvhKhQxBt2rc8CLg9p41MYovMpx08kZXLCsGHOYhiR6et48rzbaJPumaCEi3qcxsP
On5kRc0yEYo8WUcGHuOaNqkuhBeIDZlyOhjaGQ2NdM3jAi4k3BvADkjzQ1m2zucQEsh83UDlf7GH
b0RE1xGlT7el8tXPK2yVogaRCQFRSEctsfy2abCia35WKlTQiVgLAq/TGxLi30cTRQUikJ92PliS
wjQ98AawVD+g3qC+GDR5gvYesH8YhF1B1lMllCAx5ZPYBsqHkxRYA5uJu5agLANT2rq4LEdt78Da
Jtstm8WpZxT0A5PYEHYfjiKmy5eqZKYcfziROOTbCYWQIskwlejd/2tvdPN9XdHu7YHNgYsuDJRc
oHUb6tlOzwkhl0VJWGx7Fkoqy5uIMnv0tWljNW7zgOFo7F/CIHAkFX7l2cZekE5Faz4Ky2qlSIOB
OiRb/+Mmr3gQ9nOnsL6YhlpSXn1Bc2N6xkCuSabSYLzT1oGTY5SI9RpAaB4xM7ojS8+G3vKcTyWs
NTKKC9jrgoMxQfQEKyjNx23iH8FnYCNgCl69LPA6c0hSxM1174CuT6QYxPCGUBdv24V7uK51n78/
Scteoa64pGTO05pB26GAn5yLTZRLbxibOxsFSVJLVbJ39eNckkxDgnpZD9iZ6MjyDusmu9bRsmiA
b7gtsEcwlE3Te/nO1SZcvQs8pGzEUeFG9C9FqT/rOOg2/tKlI+OlOgkz1qh/9h/4ewqp/HD5uOWF
lvamSNeVw3GitK67ly8E5MvI2K2NU/cJANBI/WIXk64yXeCzD9D/UiNA7rp04vpVVDN0ggwHHBLg
SPrzeQs/wQq1lZrwSuZ9NDniyKN12sK4td/5DkYilZmgzqTi2/mvkLfE/+xGulZHntOLJoOyQQA7
XRkNz+ooKjpLcr/yAmoh2R40sXh52yulzWhb4A3FRS/KQ3wwRnrSaX+mbT+wA3rdBS/4BaXfj9qg
dXuMhBoJhefyMpooYWQD3XfVnhtjOf1U5apyEQH8B/lDHdE51OL7E/lbLTZTIx2IO5HVbXw7cSv2
04rNrL++Q1gI/fY22M3B/odaIxp/AXlqEC2B1mAjRGtbWwCvKlRKxp8MY/QkcT0fH6fsvoQUHed3
KfFidGY2s1tSBmmfGUwga/2X0of6YS8/+FPV1PQxqZUJo5VefIOV/h7p5vFOHng+pUEkKDj2d/Xl
3Rg6Dsi7a+b0FyYaej8PaAOR73E+/yQX40lxTCOlQ2Tl8eWI8SRZkEzhUQX279xCrHTHnrQGmzwI
Bg0KHaH5rdKHwKG89Lhonunh0SCPlDJSws4QUNoLFbtsL2iqC+NtjQeZHpSkOf0PHS43Zv03GfLP
iMJ/f2Jz+LvlLLGJbYp048LvfvyaSayvsrvttN6y+P5g4OFT0DM5kDaBoQcv/Bo3yHuPE+n/3Fwi
yPbs7uEvJ7ntmNZIZcDDRyahyuqYYeeGpf1Z+VopCK9T2Xz/Bzn7MCg1BUt0ME39jqu5DjbUxHax
ElNRdzpN4rnH4oJwcG3FGdHGZVvOlTaAdgQVCnQ5c4V9NGSoni/deold7S+6pQyHG3RuoJ0i/gi6
akHuQJ3t/pBjcGgA+ho992hKUm8j6M5vZfNsEk8XoidW15QO5+K8xgxP35fPQF5uZGm1V8t5rgub
kcIa07idFWaIfWWHazzViB8uaIVzWdU8/aHEKdUbMoHWXg3AfH9MmF1QF6HlcydrNQM5XVByMtF8
gJyPp9RQ55I/WEE9JqjU84DM1yQR9NUjSVYt8b+PWLN70P0M3AAu0xNr7MYByqLQs3D6YM43Q2Cc
PAp7DA9jKLgJVv8jcxUS7B1EEgk8C71r8YK5zmqBt6l7TPcyBb40bXvNhtc6dwHMCWAoDN9SbCgr
/oX/V7KQSEJWwrWD5PuVqWbN+NardNqlLe7ScHEl14hHbZpxb5MuTAnHffh+zc3yz99VWPrQxTS7
Wc0Iao0i3ph33Xj1I8NTMo1I/x7YxxrI6BPtTllLdcZOjVdXYtBrVVTLCFWROClwpd+1ahzlFp9L
X7g/Dul3sNTHr9Gk7LthEUklT5S6mowFdwkrW488LAOvaAHh98M2/8oU+NEu+9KfTK3uzef0P86u
hLcLxKWffvgnUtqQqtGTqJsg56Wu675CJg3MWfhqP8SjXhVGTyrVCt7Ph2XR/gnRECFKDyIvIMAQ
QvkICNZCczcb/enXOPAKMmN1yMvHhL0JaLLwMH0Jt3COsI+hj6ra/M7lu3cqxcAINfD5k/mZ3tE0
9r3Attub/ZodYddDTwUmpI/L+jko/JJlbl9nplxV8C5QdHsU6p2vFInPog2jecB91itnRal1UHgl
KGdXWv3d+c1Y5GEBiXoUvnP8Ol3X844H9CXUto9ez2IM4K6kAg4n5xkMy0e/hSB2K6rMxxZaUr24
n2rDfCBKww5tIIUIDE1wAXgSjKYhlZKHB/Fh2xK51BatKvpj+nuZMZyhmxwd77O7T2xsUEjAvDWz
8IRKb+7gmb6mknrejmxbiMtYsGAQ666hURtHdhaLIfc9grKR5wjvdDYiZSTf9O9zREdjFMSIT7/w
2UBsMOOhmWs9o/QuzFLf+S2eoO9pn/fuhCTP4eIPV8NdHNy4msE67U0/rhMS2CBeOe0j84e5TJvv
4DD3/o4N7khejFEMMZK7p99afh7CmzwNG0yJoH4JJSqHdKY3vKxmRMGa+RvkcRP+Y2IX00EqvDTF
kJTo0PCDrtpBFG0qEF/5Ukd1t+/5Gj6nMVoumJYXAyGITR0u/4GcQy6nho+qqynCd114CnRdyZQi
qARpTZjEOPMkr0QUg25NtCPlsB6pVaRLYsnEdSupUvGAa321eeSGpKfNSRQfvjm/BhvsOUmJpzuR
PLcNkeXxbvfoPUiNovsGmfdaiHFyl8LfIWkMkUv5baO1oiKVaYG8Y3wlOwaef+d3SyZ9FtIa0m9D
aqpM4yLEew6zBnXYCBQIiGLVyQs6pptHDt+yDmWlaBIKt49wG3MBFGxPHfkxTaurxkvM+ABauoLo
LaQDY2WjmC1Dp6LN5Rvf388mVex74hPgSAKcDMtJTe2VppCTyCk0fhR7sZy+IIlsAJS69lvD+Fxw
RlULyPi9zx5uXC51E1IEABuNLWpdFTY2kRYT143jSss+Pq+hx5nnc51OG+5EK2rx0xKSqwhBuaJY
mY4QIIiHWtcB4uCw3YatITiV03jjiYVGgrCdOFt0EryW78CQZIbdwQJ527VBcfef751MgPfhA5H+
yZdOndk7a92HpzpTtg+r78yMx7GAvfX6pJ4feKh8+ERlnh91ZN67+uVO/CmXrL206HoNpvrZIqQz
j/lo3C9GmTcNxsnHO22AKjga45V7RJ/Y+xZCgug7t8Gaw+SHu3DFhEchY2j/PG+yTAfjWZD0s1iW
1hgE4sgLSaMUXP0VDj6NuD1tpvn6q2xHAJ6IMv/j5pVyuE7Olq5OJ8w3sRVZ2Dk2B4GuPB0Y87/a
SkbMlfbyhr3kFV+ImnUBtAfhfR/ClbHupc3FttgFyXCxK3rIuBlAhXo76pChisYsTwgzGb9PcweV
cFJFTzK6DZiR7FX3PTqUBL0CWTckzOs68VA/TschPPnCLa5iXSNs7Jm6WFumzePV/RNHhqorWv0x
0lhMy1rrYa/lFuiuLsD+LJEKWmb2E1AqDzbfCGLFIEiFeLzTJ6aQgn146WFXVPE/YghtlaPHwsgg
J2ywlOelmYbc9bINoQkEGQuP5MLoRrJ6qjloPxtXk5EgiO2eaoHaTbLJbB560G7sYalrkEt0Q/hJ
RYTaH0Zv9L3aFfHXNFfDsmcwHzBwnb57bcqInHjT4qXHLfFEeiw8rkcqKSxTDGhc6mdMsJD+upXN
zGEtpXBJEKlpSoZhIi+t3cpRKglkA/y2V/i+DXeRs/LYNFJl1/yRySjkoYJAt1C4ScvetaHZOk9I
al2NRAh5isWqP144Yb8mkNLoZgu/ocGXFHzFB3uOM1evMqElr3oQkaDJV43cFb849hRhHZu9sT/N
UspvNwUmur8OIzMha3icD1lkof31voE6vUqz7DFCagdsj26jEEYdECSV1RcMAnDPv7AufqB4UYoL
auRO/UhtkrCDOcN0ZruW+1IwG2dgXwByauCPIp+S9Yc6Lhei4kSY9/QcX3jGWD58ws8k6bYpTOTk
6duntVMnZnx3QDdv4SUj1kAH2wNm7YadJ538wkDZhq/SWU9qVOUms3FZ3iVu4vyfHrsDZNENfr5P
v0lQjctFq2lkBiPtHyXdSHzuBGeGgdDYaBT2do4H3R3HY7QYCj4c1sf5cCVMbr3uhIyhVinukEOk
etMSqTVrJkdLK/yiJPqM/GwHuYkf0/dDNO6SRCBNXaiGxvQ1OTbMH03kUCZ7BvlsKUd1W2sxjC9s
V3+g9UBdEnG4PU6m5IoPqpB+7YVxfXY71wtJ/yPphv+8g89z5ARPJDdsE64PQ1LUQky2AvYTzQeD
3pfDO7N+4bSp9n6lx//xRT8mwQyMy6G/zYN5Xa8F8U60/D9tg9HedZofI70dop+Gc4MeTwvnhsPO
rvxAeX1jBowB1leIR1KKo4G0344bpJeDt8+btI7M55USk6QFisWE94joHiCXEZh/5uWF8i59/hgj
svC03ginGHh11EJX5Iei25Yu9Jj4vOSom9OqYyu90Ka/AFUsD9R4NTmZMa2T4BVraGu19uCPkIuD
Xk54/75wvwpPKqpXIrjtbycgVvB14wW9hQbe7YuHU/Re5Rl959addctsdnzTU9T9+FjGkQT4QYKX
i/XHF2dT1Ry+yNx37QASD2lwdRLuwE3UeFvTlB6Z5/Nc3c8lMRQmooCdfy5NxGCTunEaj9dqCQod
sGCWu1VT+6Bg77DmdmtdsIj0EPA+8AWvdCBLXamnGTHMDSHNWpzzlU+8kKKrAljbtnNoLj2/VNUB
2RVmqJvQANsjSXUL2s1SLAGxVuGtG6OW9IaTMRCVPbY/Ezcx0/6qBIdCafasliFebYPuW/uiHlC5
C4Bz85f9yjPs1+WPVM0QgZnJXBbMKYqpc11A27ReuFD6CK/Dyp8YTHQIlrkLIC1qjG72qY8EZcLf
E0RJrjE/WR/rXTOh059GjIFNJh7sQeJgQbBJGoJi79WqSvLWrhdX4IYQEKAe4uZP4Io2fT56utYk
Sh90HvzgZ0kz5iL6q0VIK55ItbZZUIrz7izYFKJvXaWGFz481vL7/frtc7w4v/9HdH9mFEB6vn1f
m9TBhjv4bB1cbqQTbAyMkazubJHvOlsdmJl5AX0dByt7Odi4Ek2HhC7LxbyTOJo/GA5dqLT2nnY8
QE8Lit2vTjyMmfrWpjswDn6IBWv1EDsyL6pO70VJHsZhHWdWmDJZuH7/yrdbDTJFNalMrTIFchNA
4jBFdodCtSPj4YdX5Tv3mCsv5upwp07SV4bO68aTv68vEFi8JC5tKcYB21ZkRQq/lao4aV2Us+/j
94o4BXp6BG2EiO/95kqqH6jdghLfSyi3CAzzp7raCR6dRC25KoBoNcSbg5FdaBBG/Y0hUdBfRFr2
xLMQ+dH8dZ07M5iEc1IQB/ojc48Vkwdt/20+auy4dcer747aHD8XvGSD8vStUCbdqu5JeH4BhR5i
3L97qRoUG2KFXpw06SqNKz0s1vaM7RfD4RcsD0ip2pXLfgseuX+RKX+mSUmtgpBKyC6o7epHbZSE
GM2gar+Ir32+dXUhPToBU4EEVA21bLPlcjEzYLkGETRQRxBMVH/isQ4mrIDMWXK19V9LbPc3/l70
EMCEF6lUvIDdLRQkNqmm7mqK0ldhi1PlJXTcGcDDcsGC7Hnyyp9uFtRvnyZ/oIWe/AGH3c1K/W6D
bKqXjdcNQn9/DVoK4Npf9kEWlHHm7xcGQ3nxNiWIHDMPBOIv9D7Mx/jl1i6iAZYhAbiHCWS7KEVI
y3e5StiPYp/TMdGeIP90IM6oGy6LZte2ctL/lvs+YKjbEa1FAZHziD7bWc8wTAWJlj/KehJnxov4
2VFvxPRhVNb0z9G2ymFlVcjRozTOo8L+RlBt9RmELqzTLdifXNRhg6Q/857psxkOwGYXD3QXhlVv
yx2fDSmuxDThQeKvi4AZp1G0wor7Bon5ECs26torA0rmQG6osK5kLhtGcvsNyd1JVjp8sCj1T09/
ReUqfXdlEMt26gxbr0adZW5uenqgbxQlcLU73fo6/KdaIiXqyqBgB7Cie6N5hBqNF0Fl0lN+NKtf
xluMJIBbWEHCX3y8+gJYu0qk8f3jHLrQ0gTzWsDwmLhn9HS4iZlXzVwW/EPH98DyXg8IX+VE7tWk
mq02DP56K0pWiHQ0JS1QwCNhc7ZoCV2dlgiEGNTalcUSWr2h3CFntacR7tuFWxlm++YXGDATY8MU
CNUvGGGN9dc7zilPzYy3znKqGGBIrOExKfvDqWs8h5+L5Zhbv8sEA+LWZY33ThDl0+r2Qcf6CPxo
By2DTsEflfd5FNlOd1jLC2cFkCiAYL13YYbII9Ne6qsPBlaoa7cRuuy/1MsoVtdVSa6hJDBrHOF/
+Xthp3lSBJbDATHsGEP1VLsGO7yI6FKry1nr/uErGXhV/aYZC7WeCpTFsEqtq5FtHoM0k6AsNWz1
Z92JGGGHTMqPY+/bEfBWRkKDQQl4k+Dr/SzyjiD9J8tGSdEfy+Ekx5zH2oYJ9cfpIuqKDUoMw1jT
1WCLle4WmqZZPaiD4DFli/ya+YMb5Tnx8X41Ei2nvsdJieGvSJUC3DwE9edx9Q9GooyqvSRdBU9S
k6gbxS9sJD8v2UztBMJs/N84a74Kph3d1HzF+ei1OIfkmlohy7qlMDf7qIc/HrCI98McCPx6TF+d
tLHjaCFZZQ5YcHcDIluT45/ZsRjrKHJeeDzQc/DCLVED8SOBDKHo8Kk37BkROI4dmPVM/roLNPXr
I3YTaEWWvhgZZ0iSZIjPs9h/8t904bO4MMYv8YsoPS8ENp9O4SXsPHWJg7ieipaFXr3IxzF0L1WA
ksu+cAFvkjw0mbVb8mB/IhvXgzLiNuAGGHBHFDSDgx0EA8FjKruh/IU0mS0elWgI2T5ogrIFGHgY
8a0sVsSPFvDAct1I8hJ4/CUtb7bio0fLAaa0c4h0aZpP73KpEPYktM7yzhs7sZum0RrZzIwt5OGq
LxtGJ1y0M+hHH58vb0WGBjSkboMSwvz7Xt5U0Yk4seAb19ony6KOrZHvnx5S5E/ZGldO0muf7ctl
8pnwKGl7TanrJ0nKxz/VRs4vflFlbObzUY6Snmt3A+ghg46nCp61tWwucRsRxhi/5mJBIQemc/qM
273lBRRkZ2OtmNDYh3iaEsusQFXcx9NEDSGHT8oAZA8V3Kd4aTocJMIpzrI4I/Kd9oA/rtgVfIT0
2BIaCIcpYzelNJiJRPiTYZTn+eTt1tNCC/aaPQvhcnuZp3RA35SPDST8rEisY+Lj04Bw7DGPDx13
Hk43m5ZT+nfJfiREjHlKL71ZMDyLwAhdMp4kDIg/sIy+6gW79qyKq9bVNGUfVVLDLniMDbChY9kg
UkacsZDZjdbTJU9u0K/+0NL4z/w+VWaRDCVBBgmJcik/CDf6gdJHP8Dufltm1DfyEC7bwqrgo83F
0FhMqNX0UIQCr7kEcPpCCwKMl5HLBGttxe19cstE+QpElfgvLvaG9no5zG5R8OZW5L1XXeKuL9U/
JVxxM47XxdNmNA57EtgNpNms2MdfwLIQBe4MTeHMiFVPFP120/4q86PD/cVpFa+/A//OIhFoUE49
QXPxLrdyLnwOSsQ7bxNNFIkKmAH1tBuzpw7Qz114QuxhnuUYs1M25rCMRIcpKpld6cOg5cliwVjr
/v5HqP7awENYBS6W17Qk+psb2fbqV6TnL7CDaPnMeNY8aDa5pqVGDrb7EL7C56OqWTggwJqPvCH5
gtMeJ5CZ5cbwaGoDl8okEs8kwePoftMHHAGgsZ/mG6glUdWBo3EYtQ1ry8tLg7yy/QTstXscIx9K
+fv8BKlMaY0fEas8/Kv6KzpeQvHdgX6rUrLko+k4H0oEMtXqqrtLhEBjt4Z4TreSLdVcMPZZbd61
tRhFUATkCuKRFC/iTkC3uBFzf0Kjoa/vKaopj4VZs5o+MUXinQ8b9wHYKPQa4nBw5JI78z7O1X0Y
IGot+MhRrgVKucBkyef+JoGU5G/EuQlpVtBzv0YVSrYOy1OrZl5KtICco91bXkKwDHjYmbcVgfaU
yW/W4YRj9g/QBFbsNW7CNWkt1PozZM8U6AQFPIvw9AXMnq1YsCZZwkboyvhT5nnRrFISvNWMVw5P
0EafEJXAx5V+A05JoqXLze1VbKuRMR9RUrqqvaSMBfFPCm4Tv5pnyO65S04rPOUt6xzSkhQKK8WN
81VRLVNvqrYsqsNiCWJcP7+9VV9Fs5E0mEbUXJW/6Uoj1u0VqrO2jXZHmNOcNjFV6iEtQxZ+G3jd
ttgDaMfr4WGvJ4q52kMRZo8Ni1AuLROD09gwsIGjxLqLfzEuUzkkCnV+sms4zoHf4+vX6VlZWa92
pX0Zg49B71KYXGkmdDsLZPnpZgF6hMFPLT/wQpH51dSZAzlqj9C15fT0WvpjXvL0+CuSGmv00QLt
XY78PJGu5urFcCCoAOgM1ymz95h6RMFPAlWCL2AeOg34Z+crECePlt6/0EX0cVKg4poTnbdlspl8
m6eC54E+IuMBA7pRmXyBOaQ9pYSy0zzigSPr04oOqiroRrgcAOZdZCMxW6yiLV+4dDEpkR6LT5By
nVVSlD9rAkX7MejwWKdppKshqX5vKKH6nIIR6C3w0GbKwXgZl3nE60PkcWdlkDjLYjHRp6knkqWs
h3A4us69LNOSDkL2tuGh89MunFAt86YZTDNVScxFJLyYsdB+msF9Jug1/frqdzO7VTOqk32T4jaC
CVYVyx/b4FbfKhjAd10MAENzC/hyTzvSqhfZVhGVrJtaJCnFNoiwLdfgpk9mnn3MZnfXpgtXCtuv
cr4z40rQz4fJLN7VDCsgYYY3Y8qvQ20SKgQyYfqEMGyw3Z1OugbHAZidZGeun2n3N/0hk0dsREyd
eqXW8ie3+Qzpi/XR9UxrJUXZ1WKGgC3O1GxnQ7vIu9kOFpUE9TrbDiWRMORSbm0tSF2AbluhFjME
GAloFbAX9IX5uqLp3yZEwCtiGF/HvTlEYMXsXH+5N5o1t0tLWbG1P2vOPvuhL5z+DlOHtYqllOC3
Vl3MnWDH+sS3fbwxyT5WENQ+RINBcQOoRGlT3flEwtVIoAj2Utg98fmsG3Hib8G5UYrGEVFq141y
OvUzylpDPvwuZdb+LKknlleL1CryWvuYvIJCJl6zbZtVzru7n+oTisi8X8SqZS2sqLSkAevtNyUV
LpIjYuMgezgOnX2Gi7Y0rswtFEVfbRpNGsvljBsv2NSermqHiTIrMHjisKViaEVWXPr4dSVDh01L
GVVdhUqYPlYDBsUE0Lp4i+EJM524UADNgj6Z9WxGcUYIjMDMYC9WaEzxD+u45StL+IWJj7p6904x
h6lScDBVwL7xvSdH8jber1ZuWsPM7i04Y0zqC4r1gNFQIc/LbR9UM9qlxxa7LVfjLKZRkvzMxVDb
cMuA6whqgUv/Y7W8T1uZA7BfR3Vrq7Rw7U5chmMfXiyz/8BCr/7biC27uFQhPIfW7UzCAbpNBkA5
7l8UkaFiLVpVDKnDuWyvFSYxzinSJSJcOkgIYpMA1/HK0cZqAHDJiwZHgYe/ySr6Wb/NOIB77UKs
BdAiYQXoKk0P08rT5SV6I3+tHDN9QeJ9p1j6jG2QaSVwe/jNTdwi05Vxv1XlSNLTjAS9+5Ctm+F2
pOpDhVg7Vvxc+BIdOKV/QJ8pXD4DSgar+uBiWi/3N5dlbGb6P/BeJ+FBjC/8+U9Xe7KybduteD50
X/PefgDV3teph6vKrQg0vJk1ebkUy+7VnE6LYFCINju9Bj225xIBRFICaeoca14W0sqrsgXqFcGf
CCQ8Qg1Z5U5KGlE63/cw2zCKBeEGiDftoT3+2R2340odrB5EmcRvutniNOsW4yeRzqPgfAuA0xSG
WhtbpA9/kxf6Ta5ntOkPgNmdwu8wHOwC5UxwB57xJ2rmhNeQFsihyobRe4rqjCudNHahhfHOFg8V
JzdN95apHwgG0mtl5yQ7U5lmoozzHpq5TzfHOiG7hO33Xqv12KxVHgg2QaWyML9HUmyM0pv6YN0P
Go8E+4/W2MbqodxL1yzThcC+0B07r+G3TfCpU2Lm2OPQHMgjtpBMIwiVD0Lt4xGK0H3Q0lOTtfQd
Kv3066wvNjmLHepy7rA+Jf/swaPfz5xN1M+RMeK/LRqmnh5HL6/7Yj0u3NK8A0I3A+yQBaz6EOMn
YoBnC0k2JAEJ3C9NtsIqLGLaVfvJ6aLdtsNKCSEoH+2JzxxN0HHa2RcZBVc+5Nb0oXagvteNJAz5
0CzkazML5tkihP7ecH836wK56z6x+ljFGKyIs0336PEk3y6jB6qO20ILvsCOb7+7NhemvsFMOYye
mY+A2qM7FMx/K9c7e33bJFxeBWg3efNlpFVyXhk/Q/Vl4zysCsj/BdIFch/QkkxIfx3NOMaz0vPd
QHdY3+cMWFLj5RrvNq8h+2bMViLEvV7hAxW6v0Tk/qwUdNLk0UZ/tQUFLKw3dTDHstOYwg/6Pupc
cB2oglbp59xT5sqHoBZgjvkg5ed2ImOAbiMr5FU+RBL3J9gcQNyjMJKAVpDeFp8LwpFwxNaYpxHb
q4fD7hdtlLTCTh1fdoKKfasxHeh1gxssSe+kM4HPCNXn5HZpt11vkKVHOSdjyVCUTXmxWU4uQkxa
DNJwhQm9LgIm/xs5XUMXgXnz3T2c1j0482K6yTcWjj0y0eqQt7IoFBn94kBrAZvE5f11dZExG47/
pvlHjFbLO+E4Qy5DUBmxqBbMn0FgVwUl7g5iBoCZEcXVXNW3jX5G83uplFOeKepeDUOhyptgvBue
P+vbNRgwhFvdQvQRbiuA9ReMjJIw94YkexNF+8V81XD9OlS7PFKCfAd8DpYIfsNHhzbOywlScBwq
Rir8j9Yi89eqGacB/+cld0sn5/hbxF7gp6bR7pAgr/SPkOj7bMZi1QTWuVv0bKFb38L/M/DUreld
xp2ptlYybHHFTifQC9NAg4bkJRUMDMuz9kxWdCdQ7LwPF23z+w+dk5hEoF2Vhg51Ha+1vyMfmbC+
lbB3N11pSkIqmBwOFXGQFiDTLBn0fkaKUWdNE2+0/b8+OBY6g0i6/l9B7YnsHXK+6c42m1ttQQ9c
wBxUr5vvFRnejhYDabkKT56sWXauPgs0vCGEEovuOT0OOPXnRTdtc7oLQYZFS95Q3erOOzcj+Pqn
Wkl9lj3096/3HdziWGntxLSi7HR427peChs5i4moHNNhlQUMS8sPdZd9OtuxVAPmzq54IO4W00Vc
6t+aAw4LfsmalKHXSAIDpkIHT+Eg3eYR8fvFBrYp3TR+3nrMYoeRdTgsdfpddfB9oE440P41liCZ
VoIIL2WNoCUnjdRp2PAWANzZcJNPUnD9v9kHXX6J5sBMFnqyVSrk+cMf6jMKRGj7fCF+bu9g9QA9
ejTNK5n/sYsh52mX6BF0RWTanrobMPYljhNzxeiSqx+T+Hi8ner+EI8rYGDNaX11Vfc5bCrjvpGd
HWmK8XEw+m743SUBx91nmHeMrw1YQsdgBhdjpDRnP049MAuS1bK0nXQj5Ua+VlLP18eQXhwlb/MH
xYHJYW4vNZAn+NdUvsvL3UAS4g0GAGo+047MY+F6CyNBvg3IE7T34uVzoJ/60qbiIVeZ6zrKsQjT
bHrmxjktGMMGh5itEsDXYQ/We//v6eQqmWjsBfaugWIRyQPoFL4zUCHTRymPuAjH3DVluWsdGZBs
U9g1MCX+bXihYAaWpgcpb3u29VI7MTaTiCcf0FKjbHSN98wi8M96ofmhdP2KP8PhkKS3iXbrNsij
tojJicPznSNNnwf04u/zEJqotdZpx06YFF3AVXp2M2+Ap6Ig1q8t28ZxK1ct3Z3akD6TVM+OX30F
GS4XV2qN9EY3Br3zM1O8EH4HCMU5EzKuysaIJDzFQ/MSYtdgLbHFusMr6yp8r0aKK78g1tiAiklj
ZTw+c1iP/cSXvseDQpkLEs5qGF3dKfFPj8VFklS8KNidCSypwNvL1n3h04bLbRhVFtXEaIPleUoT
Wd5fhdg0cBOeCMbmWoDgqOHAGfHbT/7w/5b3zG6alie+tRAg2Ft+b0OvHVy/Ytfxp68RxkWo76H9
zlvxYRfMMUCVz/aOL7wsm3IOaB5LaYGp7Qk4DgwOr8blSgpNBWqwmzhQ5Or7pOKxkpkUSbefcYd+
EkRifmsX1bVGWIoPgJrMBaVFiRUODPpnUJxV5cMGRyKHo1O38n6VaRbe1L9iW7WL5MpA19b2oi9B
T/QSyFdg+htv3OQl4urf3J9liuuckGpBWStxv/bkMOKeFdcRBxeCitHRtsYIxX0HWbgye6NXAS+L
yDx2tlPLC7zlXkHA8R7nBSgIe+MEQ9sjX6LBMQqif33NSff/UEpR45NlmDLmVuDL/RTuzkHIlnq9
qMacW9krGj5zV77t5r0tdW/ismPMsEFzGJERatSZPLD2eaN/Py/OV0z5IrfXmiw0VtpS6ThspTSI
ZA6QB07WebUZ0yF3zw78wl1oyTlZE0y5Gh8s0UzIYRU2jdOY7BIeQBvoR8Pyazk51Nud2vTkzLTX
7XEA+tEhqUR635UfNI7iOkkEfuwvRWXPm16g3LfZ5/kME2kI2IWx2pxy8QIIRMub3Rasincg4m4c
LTzWPDLt1+OEtU3Oyow1OUyeimRog1u/6WlLHNlEmAr+VNUwk7f5ypJbS6tyMdm5fOkSzZ4AEMPC
np9ayH1RFnXMx2dbkx6W+lrd5CaNfkEVX9bff6v2sbdwbieqpcQbZtslKcrKSEd92fOK0eLiZsdC
tUMpukM9+iixQOw6wp2lgr5BcdsR8JJv70KDrk5ya/jKYT+sTb7mVNdf5eq2t8Us7Q4B8lXDcQfW
/HDxvC1yqmFMkOn8WLIpSyGUXnWo4jwRY1MmUgThm88bINzggC2DgZgP1op7XPutV3YFJa7d2DZg
VBGEvugJEJM9niHXECzgMcFqiCYoJ20qSxGQztznQGxG3FWfUID0T+8LgUdRmVULgAq/dvJH+4Gs
MGN0yOdl4AOANoTJKYSjLo1Zgv2rh0o1LJlZ5DBnwvhzmLdKl65saLH6Sg5hi2Oxd7q0PwDCNekm
H2TxpWxicrCP6ISaidIe8xyRL7PQ6IIiz0QSCi/JPAtTe+FqXz52+4yGdeBzG9t5+zZ1DrpprTuI
PFDDtnkmgTZ0IkYgtVw62f+1oYCbm+sp+N3FHk7njn9FQpFjG2J6yRIxK7XF7ohxZcpzVLFiugNq
1TvfeMDCDi0zXEUwW8iYFCqTkgh2iK6eq32XbkHikHLehJyGkLT/RxzxWzapyl8aVUn1tvVYnW5S
gNroG1gGcNR6yKpMlW3TcrpSZtnOdShEPpOM1xpqX7kyPf+a94EWoI7AtKgi9YyFfZJMjbxta0l/
+IqJqlf/1A7EFVhqYGpC/dqvSnDLE18pBFiE4HG15QBoMBu9iMEZnbwMUgvdALwxEoNMquwyPZD7
25VGeE3OfpHlWKISAul5rJsenmcKi+or1r/Axec34QfRfRfKa2dDt8dMjcaYYXCAijtX/qyYdxUy
gCEH5rgBwU9nGyJbfUi2A2CVuOOrR2veBTGFXLeroiGgh6xjoFkTfAk64wPOaj2hVId4N43bBHNc
jHavA0R+pOtftG82pywXIuFPa41bl+UVq/KxBXjjDQTB0sxTuul4RlzHoy/ynV8TsWLutfSXUP9+
Nii2M6vlfDwKC/ZfE39mmDAvNINDeGvvhsbzLsxKoS0/I9W6e9cdNb8P6jAfeYy78RAsIiWoobWg
+8cy7xalpwbba+C3vI6jSZvIsIoi/xJoDD6KxrWvtURURG3U8LNSlFBzRceLzwpJ4+5aVshp6erC
xaE3swXoZ5po3RS1qY1GbcKYaC5Reji6vgcJ/noxXdg1vRONK+sPJjDvgGeJTcC3eFhDVgC9i17N
XLnFuXKBoeXFclHYri+lsh/Jjft89cdiCYA6bpS1Rg/eNQL1MLf1bwn4P3dt0ZautCPSJSnCreyU
ZaXfmFZfYC4v0lMEW8nVEgocV295KI3WOtpS70+t32qxI/xtXImwMvWsQ2B0HfNH/03YTV8RosTH
yXmCSfEx+jYiM4UJXC4SxUiA6zwjw2EGKS9Ym7OSPksLGAU93MYu5pAzimkSlyTSQ+mAqDeiUVYs
jQ8i6r9C4FPLt1m0cnOu90OcR+YdkUcKC+IoCoe6PItUQjlntAT7NHJKTyLTvlIb3bXGxbSMlbS8
rBHHPJHkY71xkiMCCO0oZZPWiMc8TV6J2q/3BGL9NyNBeiZCcEjcpKapnrv9feUFIvGWorecl1FU
ixqmUhBmybmCUYu1EEdiIwT2rWVN1r8fqs2wJG9mSSzG3YEUd8WVEh5pNlnY7lbQqQydA+dinJfQ
y4F/BwXF4HC4p9crz2dNehnEuzr6WnbLaW+c27tjauZ37GmgLQL1eJ18pwcpGork8vzt6sVlUcIq
KCiyHYDX8EwwcQXnWnloyxtpB8hg8JKgtDOhB0L/5EkWn9DJTSl48QSmhqiCNvYDITAIlObfKEYC
XF+kRO2AeUVvmB9GgvLSxCy6soSd9RRr2ULSngScYNXJPL9rUMd4sv0p+4CLImFtD9706F9797Jo
2sMG2nYPJ39PsHGc3vG+oQJbqUr2x1nwQF50VLdpoRcPM3oknMtMQeNxXT2omLGuG69QdLWPPkAf
FCap7Ef93oZVyUVBxYJk/kWa+h2CqaLksQH7fuA4gw8nXC1eGNzMn3+YMk1EVOBIDqc10U6afnRB
pKyTfNUZMNjUfIsCuS7w4zGEm+jupJNkPOwRENLqDgSNhoFSsZykpN2kxDlDysyVygggwyvXPmWv
2l6sq4Q+rjOgf5Q/sGM+fbXgP5R16r17nF8JvaJx4gEYHfyoVwZvq0E1Bw4f4mIiOdj1+Zgs1rMg
/OLDNtOFEG5lUlyaUJc0ZB38bZYVd4Ygs4sGyMXIfS05AuRnRIymLcDNxtnq+G0C/tg1h48w4eBf
6djVqCs0aqx0tyfgxZ1fuTQkGmeU3bwL0TPPAnmM7qI5RZEGXJwJMyZ1jMC6pO4g8Zp5vUh1HU+4
0yAI67IBfStsZXOot6BzJe+lZFanag+R6fbRzqWkNVxsOK3BAzGxMphJNjK0LMdlL2rFP1n4aR4J
CmDJ2FjctyjwXfckLOCfft8xpa6K5YOzbSFEzahet+sFsOyUitmR12X01BN8hj2JBs2x9idYCrr4
K2DGJzSkuEzuCZwh0vEGiEnecyi2WZSn752KEkJ0b5rTySmi2Via3J0JsqbAW4rSXtvag7bHUw4T
cAeWbSk35WOWbkjfelOjBgyp59e21mLTKNiOokRIpCVJI/ysSkFdYX0gMoQ3fWNoZ65MZpp13k0W
fBIvAC9nabYgh6NG3F7uKzECnIYDhWSjoXRP7tG3PE2eg22ttAAi4QPWZqgzxm/tE79L+vatnOwV
YnKby4bSBfJX0bm8avwL3dcwwDjQMvzVxmo5YBKyuuy7y5oPgCKtGS50Eae9hemFfh1ESUwwbFzJ
EkiGwoSwlEFnl7aet5Ne/HMnALb7WFop8m1+d8LwX29Wg+T3H1X4sdeZjNliBIuxSA0LRtzQorlQ
q9VKkjMbhTIIvp1p7561h51SVZ6Doc1ykIHjdKxjWVxFPXsefWJF3QdJ+4Us4Un7VeO/d17RMESe
HFllx5P3Kqu3DooYLYyRvSq8/xc3ApxOx+ySQZ1gz5QVv5FDUqSm3BZW1xjLulikS1WKaY9Xv3AJ
+BHKJeqn4EHGTOHF6FmnNWHQ88ZwCkUbmkUFE77Ky48yShG/guf1IpqHzk65eZL1NVJSs/a93BFr
ivNYVSX67Ejjy6iwCt7eU5j4+gtJ6cIgItCHYsnuQlZdFnO3lGcelSea64D/VCBQXm3Von3DwoL7
pz1MUf95jim0eIIASQ2LFVhd7cy1ypM5pU5Q1kqArFbMH70Obp0aUM5hcFerjA7TY1qi0OQ7hrEK
POn5Llx7V32enwxgO/Z+h5+aCYST2sopRTqE7MD9VeqJ82spA81UMpwSj/h1MHo+900bywjShigv
Yj4AYulSHabpp354lkxDoYUAM4Ee8+XJwMzloxJe7Ye99IX4TvsNNRJJSTblqvweHkFintI5/HdI
7o8ggGMlQGihGn9ggb/NZJ7Zt5IzbTK2KpE4moNh3HphnM+bE+3n3JIPlpY+gA7wGpztqRJjfz4h
fx6n6No2hl+ylMgqnjbl5vnG41Uh/OgOPPQRjAKmR9802RyvFZjfCgyGXM7k37XHj/6r3WLdSfH1
7vMZsQ/RgKa6AmcffWWoMD6BvHhJnOVXnp9zGJ5n+ZzF4jCaTW6F3vJWp3Su+KSQv21yaww3XvgR
wKidpaSF1pxbDqIlsKKC7PRB1q3rvnkHfRBtjzKtNB9thIZ6/f/bdR7Ij7Us0v2PGBMAeQyLfecY
KAcIV1ocPj/qAxP8bxiRvxSPNMB/T3gEXez++XUItigOkoxQ7sS45BL999X/nge+lCuxNfJrkE8B
N+iamtAa5JuC+HuMz5j7KcG9X3wKOxRwojd8q6LmZBOPO/Wi0lxvo7lTNzsQcWsQ/KifH78kCE36
mBImAn/Ckt65+Yk2MECfXysRv8sisgpAsVezzx0qD9m9G+dG0N+x9afsE+53i9PbBuO2XfuTKSHw
4G/uzXZLj8id6/FfIpKOHPBEuXf+5Dxdf15c/U8dg1HuPM7rP7h6OLl4asKCeD2QwnsxZoIWVWh2
+YME1A26eCmv4CQQATnV44n0PHFCRtvgEAULAn15qiNEopBY1V0gM+N2OMSm1hX/lIwvwJ8R+1Iu
nxXFx8edr46bdZymLPkolT7+jNUfHksuuCRGZhS08YohbDdhpxMnNaSz4+xf1B388+jEGWcryi9W
h025NB57iNbtjp0s2BDRMpG/euxhvtLIvJg/mtMbpHkXAzl0+GBFxlb6fzzvQDMtn6fZ1jEyYpET
V2PYqIIre9jiFktZ7yeM2j3bsZwVdxcu4pIn5X/DhoPe/ASIgPVmT9yN3ruB00bBMS6Aa1C58OsE
1AIAZNaiEtomo2Sy5GyIY7Cw+8VlvQGwge2G+a3GzANPcM8U7yJN+6quljO9bVE0qY9EvJMhzPeJ
fCBGWe7NsVlVvjsBi08s3zXd04WBuUYbCpquZM8oxTdch30Wz7ZJKu3F0OJCHGygDRhjc7QhT5xZ
bmnYWErTBgxGGJYS/xANJk6uhz8KdP1IhTC3xaxVHqSEgvfxvgqW1xiI1Tei+R3pkjpNXsN7BkG4
K8ijorJhmCzW058oRUObj8Ho6X9ZFaBDO3hzRvg7q2W2aCj10hRCAPBRI+Vbx41j/ZnRTG8+jGzn
QStBBN+PGe/I0rMcPL9nOazu67Di7jtQ074CAYBLxuorHHANvN/SZbQfKQ1wwzmYtIpjWiMdkt/l
b7afnGkeKXLOYJGD9PLBedRjbFyPK5yCG/6vK3mcLkisFH0GYDXsxaHmA5+kZqI5A5tQIv6wrCQR
g/lt103k928sl/FVg204KHlOr/lJ/xZL5eUCvjAjNwONSExSYzpTNy5+2NB8aSC6yb8iOStgrqbC
U8HCUdECxAVvE59BZA967rmFOis5CAgDlb4Exh+AI6mbr3XpKdOLyCa8FU19/7MMj/rZB0OzAJ6L
7kn17QF2/VsYDUGmyGzLyNyWEnn4Ve4RU7eZRGQefItr2Zb9hbMFg7Qgdnq7yaFCnmgA5faD99Ss
GKIGmnrZ7Ec7mvWKAiba/CTHpdkDZqE6k8pNb5VRaWtJqMV23H6injD4+bIr56J5Rs9RALLCZSOz
Qe7WQDlmVGzQ7tNel28tx3ZyAAATHPlwlJidtw8s58q9VraeqMf3Xi4xQokYCRjEdb1cMqPbARR3
QyZcpReUELBG4jISFzArDZx5p2KEGcAIP8xJlDRy54ot4GuIb1fPNDK6/Muzo42M+Z/opLZlXgqN
E/qiMwPE9iSNd6d8KccUhsiHhQ6NPOoxauGeQbpWA0t3hiCg+VYRS16oAmirSyh/Y2kbFWx3hMGj
seXZZwHPkgd1Gua4I/wncI6zQ8WxPdUVPeJceSQtktL1BRwaKQiScNXSYI8mYvv0FE4rJdZEhm/O
EWtr33Fi9OtYfMXqUc/dPfegYpCotZOHdFQfldSN1kYUn21TZQCjfkDGNTl+u49fBNvuzkD2aLGM
hSdP+GKTJguK63F2CIhAccaNHoub5suVGNYiOO7kEQYxw0XaFtSm6nOiVdX4IdpGxH0+KyGDKbnv
6Q0iRS3t5XhHjZCu2pxsTy2trKYOguNCSx39Yd6jcKRgreZGh7D1QGqv9zgYzlgGwKA9kt6yb8Si
d678vBGoeu8ymho85H2+GutUNypHFhu01Wf7ieA5LV4rZEbnqsTE3KZQwvRhTp8Z++wgrRHK3gPI
rPPhdYZtlHL39ryEtBVRPjhFByXyVFDiTZCrTydaHDdJhmS4AXarEVslfFEq4/m6KJbiXZO+/Asa
5leM3XHQvoF822L/uLAozXqqCPcnWkLGHGiJDEwDhR/YzLeoTAg2kIUHj7F0nZ2VGPMB/KdGUMaw
kC64qaugy7FPFZHGTlXILWrLCdEMKXgd/xKrx5rPGilWMsXPGBrQZvs8WjXi3HJA0VWTqEpV5o9L
ppcnwnObpXKb6nA0154NAAGg+hP1VPW67DDtSOJ0bOZZr+NjFVKkmALx6hj1qTes88eGL4Qs0tyu
lYPDYzBpgYTFXUFYgl9nqkBtB+mF4n5YcxQYk6pIjrkFconXCqXZjz6GHWKW5pcZ53/LfGRgUEfg
VZA2PKlIsCHXglBikS1Nf7m7p53JHfcsmzr/qRpwaBDU2tNzBBeIIADGOfnj77y4UlP5VoNCMJyX
QlsgsC13iIflK9ubHzcSOxVeUGiBoYIhbUDJXSjBtHRraUJG+14vO1B38z5/sK4zHrQfbfDEXvws
AbefqFBRWvRvRd/e7LLtka5twqcAIJtbFOUMX8DEtgIpHJPJirt7AbyMpnCsyMkG3GfNsOAcSrZz
wE+VpUdGE/rcXkHVCm+rUOC0Usx+mloP6FYSd78cIDrFq/jww3AKQmovjfzUIFGPASoKYas1RkEs
RlJko8dyxXtvrXTIH833YRJ+WwC9iSqDkNCcKGGxW5ksicZIAvvW6F0l58sYlyKr/WPXWlKkbkQh
Co2im//chIBvVHlyNYQfsSUwbzXIU3QBnbYwXjWWzQl95kitvMzYS6ljGY5uIV3FDKDdbasFkBxR
WFN7YM150xGMY/fBEH9J7ciMuKIOG23wb4uGyRbETCf1OR/frr0vcl9weItFlJ97fy1UgAw02mMJ
5pyyF+PcpQqOooxDQTxhDpJUA0tfVsM9jtRB/CMPa/Cx8HGRxpb4FrJwnm5uEhyEPnoY2wcc0j62
a+7C6/NjoY3Q1gyKQVW1JNbzhYlta8Q7A6QtNFLOyfw/djcKD7Jdo+cMk+umY8z6KZsQMgwLHklO
hwmLuxR2pR5EhDddfHLNe/J3CR6SUfVQ0R5VEASALZGjG8R0ZJeORFyf71NC569y+zRhvZ00ybpc
i5ExuFfsoP70uhDN9NeawlQ79BTYqKiqtumHSJ/bbhBHeeA2YSXtxpeIwkYtkDIZK5mJO7kz4SRc
f+tb05OWzhGRx+UteJuLfasVARMU5hircDvO+sVh+43++HqLlX5jF36p0F6w6kuWPwKwfjHdNsfJ
Ya3evz6h2PxpG+YWAmFNVfzH9h3i9H/CYRkPF/3QM/2ZGr22rp2/qBQd3HGrjkpkLtYICRZ4KT6r
NNJR9Ci7ap0ofia5gAXcuBpHzLPqfMUwx3XY1jOEQAY805d/2vP6H8+3fogyP94EC3FcfJP4Rmt7
5a6oIw1xB/RXtt4i3phIOH7ztBoy0Ja1cBtD0l+kIUdly09ghZV24kLJeU5kUcKVbnjD9rN7qSHq
cBxB0dX0mI0HnjwVm2WdqZ++IDRQuSL0VeaxUOe3Vw0JF5q7LSIeFupZj0brQJRYMUQ3j3YlCbwa
9u/0IsDHXvw113uSkkQEjYJqfNTU63+nB+T86VBEwSHR3hZZzZgUC87LxZs8bapXSfvbCIVVOfMy
+5IBqRHw91OQocAiHI2cMuz0ADiTk+xYI+watgY1hUCtFizTl405q/sUIZsRLjTQVHKRpoAWN96D
PkuugDzIAa85wUstIIgDTq79AfJSwDzJBdzRllCLNcVrpI/RtnzUaY2Xmt5/aJfIpUQInqoJRhTH
NFXcmg2DZq1KMIt2GFneowrROcG3au7rAM5YZJfJmXFGYEhd3Cwu7LdNh4BNsaEHoikcFwIr2oDN
8I2YP5eFUhs7UKe8F2v0Zj00o0uy8KBueegT3bsleUgd4PXywPprTf1z1Ynn/OguDyaINwXf5ajv
tnOSgUEqNPqg1Q4LwOpk66mRVPraHeN1PYUGsctRmbdHcxJCCrO8I3QG49CRJK7VymCX9jPPSb2q
63vumfFrXfUBh6ZYSjH+AhMDZA8EpbX27/JH2KCJeUd3qW2NTFswr3SAYf4i4SovFqJ5W0P6k+Ta
a92ERNHcpLJNoPQ4KkOklb7zsbZyYFRRnBiEmk2qh7IoUZAQgrFf6vF0OY6uPtA0GiezKAPEAevr
tMcd4uQ/CGMooE2cbw5NjZvG4hERdp1g6SudAP2HyiW7YL8nk7CX2acFs0GTWkPQJhItxS/GI28K
WxGHoTWStOrWkymD7yYOoDs7H6y2pW/43I3i1S5qFduJR2rjhugaeNT2TcOWu3P2fL6D8mI6vLCA
yZ5wGUt8i0k0SACBEChelKTktJIiJ20Zkal0lVuv/NbBoOAE2E+FDL9aKmnVxBkQejHHhP+NzcZf
vr8lkyvk/EAUBvDxBjALZIMx355p32cuqzxkQm0yI5KD3OBXc3DuQVd3ewZWsVVI++2Oep3ec/yu
CT/Nx5lIJnXNrFsWMCQXehLiPmcEk1cvcoBxrBzWW/OBN3Xu3Fituzf3701v8CXK+tMC/GIP8KCX
jBUTfFonIyla93Ax+DTPDBQKrqM6omGzQpIvNCMYHf2b0a0wPsK3CF5mC+2aIxNoK0I2jPpfd2aI
mKxztIa4srsxrjEopk2aiFH6zXfo3YxFEwMkleg88YpbgmXhhXAuX9/R0cmCiC+j9EIrBIUHZB3C
SbxewdBiZfEdGsT1+hFh78kFNqNmxe126zOVSWCzzinSRLLlSo8Clx31sLySThNz3AGYghLsZiOD
8LtgeBPFyhT8eHYBFPLGGu1LnnupaLIzgFZmTjw3j00pbsDvQ82dr6j0e/mDwCUgulL9VV48QiQz
oFjzHkzbRzhXjF9atiKqa5CZzZLk8D6j9PQlcSgEq61TCmhq04cxaam0hzvvTEEetHDEmM7EEhUP
vhCbIn3dkRGBDJm19GyQRvVssW7NHyEjOE4HgKISG+2+ilq9NbgwVcV1qfeVk2YvwY1I/zBCM5aL
fdXhEb32ig8On2+l03CQIP+w1iZZF2exWAfDHzmtqEmpZ92l5a61MfIR0qL5Us+x5IFJYQBAK5Os
XCvBQOwb8lVnVcgks+sRRzq0h+OA/y3sxDLyt1jgH0MSOaPmGFIoLmnoXzgOGecb68iRU0xjQeJJ
G8/uf8q5P0eJjLl+7Y3BgMDLIydxLmhts+edXFqRy6sNQ9iDQANBDJhCweurW/LMPBNHShdCivpQ
sIyi+FVOQ+zon1qql76kHEWbFIttJhEGVe2ynO9fkOHBp0DxPDNkVTeeWX7qBFUSv4MxZcRYtnbw
TqYFHI1dw6Xt58wAPleeG8HTEZ7JYXFSWARO1mJSAdvuLhB7Rf92Yp8Iqd+eh+iOV0DaM2CVy/zD
zV6tA4jXAUMBDlf1rXkhk5hIeyHijIrwD3eTD5PWIg7PEDJ1DWqnUXI+2qMssG7WoTbnnzQPq8zG
pYZBVMQJzdUBxCFZYPwM6+kIBDn3RMOxAS9Ffzrun2Hs+7wze1dEvHLaf6WSHznDx9dk2IeSfz7B
NCN5oD0R3em9ZqDYBQMi0G1aRiYUTgWqJKPwJAYypZlbBTr27KXnabMQp/rTHjYoNcpmAEfZM1CP
N9RceJrgAsLq7OPKGFhJEsMrjXXv7z70AuaabZ+D5ET5ie0EfIgPPRR/vaZ0GMVi06O1nzfD/QFb
6GaTuRSurGCJTIX7gROkOKu9arHE0GqCBQ6yOmw9juPRmvJYazkBPd/WK/8vCJcKZVH7W6FirjFH
PyWlnRMf1JTTj8qGkRYUdBHyI0uvDa0jHvRnKZ8ZYRTPmDdq0B1Lp7hRzKZjbxb4hYTrxSAIMPog
tyj2z8lXiOUWjmUoseaMSY5v4Fl0Zn8HlFBTWZgGKp7B9q9S3HJPGneK+30RLH05laHVTkuxzM5G
OuzQ5LHJ07Nyc3XSljFwQDfXOXoxWJRQBa1tWoNOtYgtsGoTRtEqtgXrOosKIWYaj132vbt9SaPB
KN406AvynI3wwXNn3IM6VAq0ocnPVqBMxBvJPHzjaQwKum8bWg9lcij3mR86sCOSdyZ+hqg7e1ax
Y7vqwpPYUC29qKbuJtdq41R55aiqdat5bqUKivd7ahzIUMUrcqZi2M9AlbNbc2lVvtau4xjDKf/Q
5yWlUgCG+5UN6eD9q9R2L9VACPXFyYbxXNLUKWVqdJZAPvNUKYDtlskVBHF2ZoRN11yQUFoOfHTK
0ZBYaIPJIemJgdzfKBCcYdIO8IETB1vD6ateBouQFkeYqPzrH7VqfeLflPNATkdIJuG56y8D0tCe
ffz8Pz8VLU0KtDULZl/1tlVhZwFOs1VpO3cAmswXHZ5d9wILKFfSVOKvaThUiZR2rtcyCr9GtAgW
p3FTTHq30AWnDCeTwPjhe1k8Vl0AvoA9rzCgRXnVll3rohutsdHPGWPeRESKCHOe9Qukls4GAoAd
NjY/W1hpvj8lEjkIXh541bF3AX46ZDw+q3MhvfKOoFeSoiaHQJ4vDQB6aay6Y+lCHzvFauOeIMVx
I0i1I1cHpCTTDb+BvubNIGTvltNR8N+CqRfMUj12PUYQLPG3TCIM2svQhta4YhpMy7PpoLlvyZ1N
mT56G0xoaG2d1tnCuXwbuSyOEL6iovralL8xyoGABVvFhUi7YKgh1JEADpfCRdv4/uyPshUoP9R2
8V9FF+hhgn+kyXPOsbi55z42NcaOuwkZ7wfsH/Gzo0DXU42hg2OA4UXGsr4UH4rJbh7pKR4q/oUg
Ili8ccH7HbARPJt4N/r6kqjbmoE76RSYZkO9iE4S5eIF7JddxJcPUKbhZfmZjWfdFmSLOYh3IwJe
GK7YGkVB+xKy3VM3nZXSSof7PCCWS4nTYxgmGdPi0u7gihP+jDcG+tITACzK0UI3oZUCU23gXQvB
p5HHTZEXu9iCtx1m+CITLkUjUVgdPlZokPzLM7cEFQrKwsACui6oY0xX3uUucmS/2xpY/0qDYVg1
d0AKOc2LT9EJaZGYPMb/zOXQ8YvdCnkc6NBisY7FyILIGXVbyydqzqoFOTQQSIRNvkU6Rx3KI4ed
UZQF09xjdJcNnsMbYrlLl3wQ0WvKqfTku0Me6bTj8qyFrdl+n2FlP/G3zzcCm+VKoHFZx6oUQ9Bx
xwHlwzzAh/sT0+24Mr/EfzETKWbAgyjGtp6bTYOYiN6ZMUTNAPR5BzekkUnel6oLywoHpfsSgUt1
Ct8jzUn9L1fnro9Bhn31OIEb33dxF6LpXy9++U4rh+LPJKgUChchcOahw+5xoK6Zw5cFeK1z80o+
PkT9v8pQEbEi9XvZbCXSK2taIKOhe2CF47NkTDy2uTgZyV5N1Cz+V2cA4PrvaTs0BUsLS0HPzSc1
PBdXhXxmkCSAVKbytbRMwljCkD3hZN09bm+O26sbSreR049Iyov1GuUu3iQs7nXookmpJdgC5YEU
5JjoIWW9JkogSNrhD1pZbq4t3MLQXTNR5xW4QrFK7OdpO7JkZ580bcwya9fHJdavgOZ78UUWzrgo
FCobqaNKBSU/CKHsIZ3lsb1rLkJ2De9zbG1JmvA0DllTZk9Vc8KAWTAH6KzqbyANahGY4/fDS1Pb
G/Q2lVdlyvC5A0N4HxnLDEIhG8ElzKnIsriMCm7VvUtHII+bq2f0JuCYNdc+YV7okqgomVnBIe5x
jhIMGbF59KVihB23gaxpWhAoBly//b46gBq/BPQxPfef1p6K3oRbga2i7AQZTdR2OXJNF0FURTlZ
BT4O+42q3fdNMZs2ic1ToyvOZghLpo7whQQdBePLZ1Mu7NYDWaOxUMlx4Q9ZXhCBOm0QTGpMcdDt
95kcG2x56RswaWcus2yu8D5Rw4eW9FWs9e4dxrnNAKkHHfnZ4WnjEnhSLHA1TAjHAikcI0B/onh9
cA52OiDcuhBS8AUx6cq2KQafEzpKe8AOskHRqom/6gO5mdgirSvrS5m67ZRgwBG1KwGQJtxZGJdh
84NfoPqYanRrjty9z3m5u5t9g2X+P0ipQR0C+A/AlN9MOn+X8YtfdiiLX5iIGhNpAdJglXT8EScu
tCgusUtswbPoEezL9btHzbqo3+VGePk+jTUXfeH5otoc7TFfBQ27hDbQjc8JLXZoLf+GzArPGBZT
LfSB/2OG/05pKaYl3z5zFIkCU0LAGKS2eGgDawDOHqELyzZhgl3SHHL9z9lq+1vY99iSlTQfVzC9
8yKtDmCeiCmKFIAf2X30NtBHwquX5vgbwNXg33m9ASLvc46in/WaVuvJKDxIbeDBg9IRKT5dOQHY
UX37ZpPR+QwrLPfhmvqJx+190rSYZiftWC9fvCjxb+Z/4dZZEDZ9OoE0lSIUIl2Wd/7UVvnkhgzB
tTinhgWaDFtWSp1ufNaBkrT7rdxRsIarKLkCFlPNg1NAfnY7FDneaP1gXUWNt800wPWI0Prkx9Gr
mbUXmfEPM3Hnp68lPUGcmljGQCzW1Z7L+6GSgLcRw07OOorgan/g+6zMP05FhtmjTux1UIUQtWTq
RM0dpId+B4uhtjdu1r8C8d2/SUVzlQitADjHA3l02QNwRc8AanwHly/CHbwcSWaawqE4K/E7To0b
mrJ8efDmjjMRp2zlHleCjcpiMeWuZW3aUOwDFFxXBvF/gGg3p7XCWijb6XvNTh8a1owCbcGRd7uR
1PumTdUpn5A0bOIWECq1ahW360Cn1WW3zMv49BvpNe76OAzarUO/prDR15uxc24lQIJQ+CXCDHoe
2beHXTKPqQ2IA2a38jJ1YACAN4yzVC02bzLb7bMe42EGCujgWP4FTpcPDCSK+UuYc7xBO+uaoJZm
umYYUPNBcNNsNe8l1IE/9Yrvf+H1m4RpzzRUPdOF0ga3GuZRXemTHCNZPlV/YSo2zJVJPK9CPwLg
T3hUgpH+g1zAD6UvqdbTpTBwsD2Qt5fniy1Cq/8Zp4Ph+FLjRiOVCS00khtfV1RCSfmU6LLLqS2M
FYdsKYVDOxCMOWRNNDqxDm4UJcE2nGkCkG7VIFRfx/h9N4C693cA6rJzuonqrG603oUzcTZwNZUl
vRAlSo0D7GVpmvG3GQOGQSqHXliEdt5DZ+ozasdnAYPSkL90KxBfzjsSHeJSh7WLSQ5xEGKfdvWJ
rzLLoRqRP5tYPIaDovWNS6evwtJP0KRiY5H46bwaKLsNcfQNVocMAs+/JFuziYiEOO/YynFd0L8f
XsBv9LFWT4NEdxRIXeY9KtidFda4feZTXinsT6LZQSoGld8Ri/BYaGn+F8tey0EappMqWqvn9jdB
d8IRj5BH2BvcH0X2Vcs/m93s9MnuBPozGzT9v6qEQjNH6ARhVwy9zM2t4PRozVzhR9zg+LINvBui
MvMcmz0aWxs5rD8jYKpXeFOi2U4dWlVktKLS0Arakl/3OF5cxeSacCdOLXYCI6Rg4CadUncXN981
SJJEl1WcXjkBhdXTe/Ys/KftYQJ2NyCSp01g3BnGJGwIT0bY/8Y+Kima8c1NOKt5DLHsw/7+OIwf
KDCH8JeEDaRJRRbyNEpP+FJdAVcdOkc24QkG1VbRe1+y6yieficg505D12LoOQi4dZ9tqjkrbAFL
HhhCAQ9CoNiUfmYhP/RO4GcV2m4sYQk3CZW0UHQN/hSvojHz8aWJxktL4M1FjxuZwCooUFd3lImK
mOcmW4pkzH3jKkEDFBb9nlzIjWpHhwf8t57R+L2Z0EO3OYd82vpkO8NhTXZggGbChsxglWTBw0eM
Bx15f2U/jVpXIQrIGADZndXZSRM0DLD9Qqf/IyjiLLPCMa/wXSqOr+HACSZqmGwogYwi8QVtW1FM
1Sly5aKezhT8tl/J/ZW45IQAo+RpChYvE/EIJEcie4TLU1R6hfS4IcUPOwYG7jmJv1aAokTf8ZUh
VkQ5kCaRKFT9gzSDMV8qhL2ZXJox1JFbghzcUVdiESs6oieaMyAU+2lMzBPg8oov5j8ANMtaDRRc
NSnZTTPoBOzUAfXAbQOVNGxFqyU7fR+qD1rWLL59yJL6niJUdTZ1jX18KUd4Y4BNMlbXi3/B6I2G
USKv7TTyqHD5lcAYXuAsEcuUbASrDDkV9sFGRkHO7MrQ0nKEOfohK8xM/1ZP9Zcx79s784kh65Ul
0e3yWmo+3hzO/rJSQA/RqRmTNZIUy0KzwDg19TjMaBrNpJLtf+fk4y2A7MECQas0umkFBG/Jf/eh
aL60CzY0nRqflAU2o1wCgWrhGKANyo/Y2YfN1purUbQ+fryV2Y7F5uf4D9apBZh9pXfkVS4oEQ2i
fBZhi7jLDLMNfDyteJN+6hYkFeXSUlhPuQw99y9hRJIuyzaX7NDPVoyWgS7qfO1rvQbReITYfoTB
wPGbZ8fOH6kBrE3pSVFpMJ8yAlCA4CuA5JbevNP4pywMTjW8Ie0FJp/wO64g6KT4i4Bl+O28YatA
FCvzNPCOTanl6F2LbdbEwUjv8hqwmrFAtyAgxfW76hYaRnnZNGnwi3mzSJKhw4xZjkIUNsnDvVdA
aF1RfxfaCgQ=
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library synplify;
use synplify.components.all;
library gw1n;
use gw1n.components.all;

entity PSRAM_Memory_Interface_HS_Top is
port(
  clk :  in std_logic;
  memory_clk :  in std_logic;
  pll_lock :  in std_logic;
  rst_n :  in std_logic;
  O_psram_ck :  out std_logic_vector(1 downto 0);
  O_psram_ck_n :  out std_logic_vector(1 downto 0);
  IO_psram_dq :  inout std_logic_vector(15 downto 0);
  IO_psram_rwds :  inout std_logic_vector(1 downto 0);
  O_psram_cs_n :  out std_logic_vector(1 downto 0);
  O_psram_reset_n :  out std_logic_vector(1 downto 0);
  wr_data :  in std_logic_vector(63 downto 0);
  rd_data :  out std_logic_vector(63 downto 0);
  rd_data_valid :  out std_logic;
  addr :  in std_logic_vector(20 downto 0);
  cmd :  in std_logic;
  cmd_en :  in std_logic;
  init_calib :  out std_logic;
  clk_out :  out std_logic;
  data_mask :  in std_logic_vector(7 downto 0));
end PSRAM_Memory_Interface_HS_Top;
architecture beh of PSRAM_Memory_Interface_HS_Top is
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
  signal NN : std_logic;
  signal NN_0 : std_logic;
  signal NN_1 : std_logic;
component \~psram_top.PSRAM_Memory_Interface_HS_Top\
port(
  memory_clk: in std_logic;
  GND_0: in std_logic;
  rst_n: in std_logic;
  pll_lock: in std_logic;
  VCC_0: in std_logic;
  cmd: in std_logic;
  cmd_en: in std_logic;
  clk: in std_logic;
  wr_data : in std_logic_vector(63 downto 0);
  addr : in std_logic_vector(20 downto 0);
  data_mask : in std_logic_vector(7 downto 0);
  clk_out: out std_logic;
  rd_data_valid: out std_logic;
  init_calib: out std_logic;
  rd_data : out std_logic_vector(63 downto 0);
  O_psram_ck : out std_logic_vector(1 downto 0);
  O_psram_ck_n : out std_logic_vector(1 downto 0);
  O_psram_cs_n : out std_logic_vector(1 downto 0);
  O_psram_reset_n : out std_logic_vector(1 downto 1);
  IO_psram_dq : inout std_logic_vector(15 downto 0);
  IO_psram_rwds : inout std_logic_vector(1 downto 0));
end component;
begin
GND_s5: GND
port map (
  G => GND_0);
VCC_s4: VCC
port map (
  V => VCC_0);
GSR_40: GSR
port map (
  GSRI => VCC_0);
u_psram_top: \~psram_top.PSRAM_Memory_Interface_HS_Top\
port map(
  memory_clk => memory_clk,
  GND_0 => GND_0,
  rst_n => rst_n,
  pll_lock => pll_lock,
  VCC_0 => VCC_0,
  cmd => cmd,
  cmd_en => cmd_en,
  clk => clk,
  wr_data(63 downto 0) => wr_data(63 downto 0),
  addr(20 downto 0) => addr(20 downto 0),
  data_mask(7 downto 0) => data_mask(7 downto 0),
  clk_out => NN_0,
  rd_data_valid => rd_data_valid,
  init_calib => NN_1,
  rd_data(63 downto 0) => rd_data(63 downto 0),
  O_psram_ck(1 downto 0) => O_psram_ck(1 downto 0),
  O_psram_ck_n(1 downto 0) => O_psram_ck_n(1 downto 0),
  O_psram_cs_n(1 downto 0) => O_psram_cs_n(1 downto 0),
  O_psram_reset_n(1) => NN,
  IO_psram_dq(15 downto 0) => IO_psram_dq(15 downto 0),
  IO_psram_rwds(1 downto 0) => IO_psram_rwds(1 downto 0));
  O_psram_reset_n(0) <= NN;
  O_psram_reset_n(1) <= NN;
  clk_out <= NN_0;
  init_calib <= NN_1;
end beh;
