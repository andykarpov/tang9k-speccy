--Copyright (C)2014-2022 Gowin Semiconductor Corporation.
--All rights reserved.
--File Title: IP file
--GOWIN Version: V1.9.8.05
--Part Number: GW1NR-LV9QN88PC6/I5
--Device: GW1NR-9C
--Created Time: Tue May 16 19:42:30 2023

library IEEE;
use IEEE.std_logic_1164.all;

entity Gowin_pROM_font is
    port (
        dout: out std_logic_vector(7 downto 0);
        clk: in std_logic;
        oce: in std_logic;
        ce: in std_logic;
        reset: in std_logic;
        ad: in std_logic_vector(10 downto 0)
    );
end Gowin_pROM_font;

architecture Behavioral of Gowin_pROM_font is

    signal prom_inst_0_dout_w: std_logic_vector(23 downto 0);
    signal gw_gnd: std_logic;
    signal prom_inst_0_AD_i: std_logic_vector(13 downto 0);
    signal prom_inst_0_DO_o: std_logic_vector(31 downto 0);

    --component declaration
    component pROM
        generic (
            READ_MODE: in bit :='0';
            BIT_WIDTH: in integer := 9;
            RESET_MODE: in string := "SYNC";
            INIT_RAM_00: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_01: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_02: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_03: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_04: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_05: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_06: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_07: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_08: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_09: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_10: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_11: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_12: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_13: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_14: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_15: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_16: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_17: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_18: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_19: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_20: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_21: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_22: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_23: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_24: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_25: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_26: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_27: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_28: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_29: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_30: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_31: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_32: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_33: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_34: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_35: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_36: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_37: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_38: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_39: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
        );
        port (
            DO: out std_logic_vector(31 downto 0);
            CLK: in std_logic;
            OCE: in std_logic;
            CE: in std_logic;
            RESET: in std_logic;
            AD: in std_logic_vector(13 downto 0)
        );
    end component;

begin
    gw_gnd <= '0';

    prom_inst_0_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    dout(7 downto 0) <= prom_inst_0_DO_o(7 downto 0) ;
    prom_inst_0_dout_w(23 downto 0) <= prom_inst_0_DO_o(31 downto 8) ;

    prom_inst_0: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 8,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"0010387CFEFEFE6C7EFFE7DBFFDBFF7E7E8199A581A5817E0000000000000000",
            INIT_RAM_01 => X"0000183C3C1800007C387CFE7C3810107C387CFEFE387C380010387CFE7C3810",
            INIT_RAM_02 => X"78CCCCCC7D0F070FFFC399BDBD99C3FF003C664242663C00FFFFE7C3C3E7FFFF",
            INIT_RAM_03 => X"995A3CE7E73C5A99C0E66763637F637FE0F07030303F333F187E183C6666663C",
            INIT_RAM_04 => X"0066006666666666183C7E18187E3C1800020E3EFE3E0E020080E0F8FEF8E080",
            INIT_RAM_05 => X"FF183C7E187E3C18007E7E7E0000000078CC386C6C38663C001B1B1B7BDBDB7F",
            INIT_RAM_06 => X"00003060FE6030000000180CFE0C180000183C7E1818181800181818187E3C18",
            INIT_RAM_07 => X"0000183C7EFFFF000000FFFF7E3C180000002466FF6624000000FEC0C0C00000",
            INIT_RAM_08 => X"00227F22227F2200000000000048240000100010101010000000000000000000",
            INIT_RAM_09 => X"0000000000201000003A442A102810000043231008646200107F117F487E0800",
            INIT_RAM_0A => X"000010107C1010000014083E0814000000080404040408000008101010100800",
            INIT_RAM_0B => X"004020100804020000100000000000000000007E000000002010100000000000",
            INIT_RAM_0C => X"003E41010E413E00007F403E01413E00007F080808180800003E61514D433E00",
            INIT_RAM_0D => X"0008080804027F00003E41417E403E00003E41017E407F0000027F4222120A00",
            INIT_RAM_0E => X"10080800000800000008000008000000003E013F41413E00003E41413E413E00",
            INIT_RAM_0F => X"0008000E01413E00002010081020000000007E007E0000000004081008040000",
            INIT_RAM_10 => X"003E414040413E00007E41417E417E0000417F4141413E00007E405E5E427E00",
            INIT_RAM_11 => X"003E414F40413E00004040407E403F00003F40407E403F00007E414141417E00",
            INIT_RAM_12 => X"0041424478444200003E410101013F00007F080808087F00004141417F414100",
            INIT_RAM_13 => X"003E414141413E0000434549516141000041414955634100003F404040404000",
            INIT_RAM_14 => X"003E41013E403E0000417E4141417E00003D424541413E0000407E4141417E00",
            INIT_RAM_15 => X"00364949414141000008142241414100003E4141414141000008080808087F00",
            INIT_RAM_16 => X"003C202020203C00007F403806017F00003E013F41414100004141413E414100",
            INIT_RAM_17 => X"00FF0000000000000000000022140800003C040404043C000002040810204000",
            INIT_RAM_18 => X"003E4140413E0000007E41417E404000003F413F013E0000007F202078211E00",
            INIT_RAM_19 => X"3E013F41413F0000002020203C201E00003E407F413E0000003F41413F010100",
            INIT_RAM_1A => X"0041427C424100003E41010101000100003E080818000800004141417E404000",
            INIT_RAM_1B => X"003E4141413E000000414141417E000000494949497E0000003E080808081800",
            INIT_RAM_1C => X"007E013E403E000000404040403E000001013F41413F000040407E41417E0000",
            INIT_RAM_1D => X"00364949414100000008142241410000003E414141410000000E1010103C1000",
            INIT_RAM_1E => X"0408083008080400007F403E017F00003E013F41414100000041413E41410000",
            INIT_RAM_1F => X"000000000814220000000000004824002010100C101020000808080008080800",
            INIT_RAM_20 => X"0040404040403F00007E41417E417E00007E41417E407F0000417F4141413E00",
            INIT_RAM_21 => X"003E41010E413E0000492A1C1C2A4900003F40407E403F0081FF414141413E00",
            INIT_RAM_22 => X"0041211109050300004142447844420000615149454349040061514945434100",
            INIT_RAM_23 => X"0041414141417F00003E414141413E00004141417F4141000041414955634100",
            INIT_RAM_24 => X"003E013F414141000008080808087F00003E414040413E0000407E4141417E00",
            INIT_RAM_25 => X"00013F4141414100033E414141414100004141413E41410000083E4949493E00",
            INIT_RAM_26 => X"0079454579414100007E41417E40C000033E494941414100003E494941414100",
            INIT_RAM_27 => X"00413F4141413F00004E515171514E00003E41010F413E00007E41417E404000",
            INIT_RAM_28 => X"00404040407F0000007E41417E443800007E41417E403800003F413F013E0000",
            INIT_RAM_29 => X"007E0106010E000000492A1C2A490000003E407F413E0000417F2222221E0000",
            INIT_RAM_2A => X"00414141211F00000041427C42410000003F414141490400003F414141410000",
            INIT_RAM_2B => X"00414141417F0000003E4141413E00000041417F414100000041414955630000",
            INIT_RAM_2C => X"FCFC000000000000FFFF000000000000FCFC0000FCFC0000FFFFC0C0C0C00000",
            INIT_RAM_2D => X"FCFC000000000000FFFFC0C0C0C00000FCFC000000000000FFFF000000000000",
            INIT_RAM_2E => X"FCFC000000000000FFFF000000000000FCFC000000000000FFFF000000000000",
            INIT_RAM_2F => X"00404040407E02000040404040407F01FCFC000000000000FFFF000000000000",
            INIT_RAM_30 => X"FCFC0C0CFCFC0C0CFFFFC0C0FFFF00000C0C0C0C0C0C0C0CC0C0C0C0C0C0C0C0",
            INIT_RAM_31 => X"FCFC0C0C0C0C0C0CFFFFC0C0C0C0C0C00000000000000000C0C0C0C0C0C0C0C0",
            INIT_RAM_32 => X"00000000FCFC0C0CC0C0C0C0FFFFC0C0FCFC0C0CFCFC0000FFFF0000FFFFC0C0",
            INIT_RAM_33 => X"003E080818001400007F080808180014FCFC0C0C0C0C0C0CFFFFC0C0C0C0C0C0",
            INIT_RAM_34 => X"000000003F36363636363636FF00000018181818FF00FF0000000000FF363636",
            INIT_RAM_35 => X"36363636FF363636363636363F000000181818181F181F00000000001F181F18",
            INIT_RAM_36 => X"FFFFFFFFFFFFFFFF181818181F00000000000000F818181818181818FF18FF18",
            INIT_RAM_37 => X"003E4178413E0000003E414078413E00F0F0F0F0F0F0F0F0FFFFFFFFFF000000",
            INIT_RAM_38 => X"3E013F414141000000080808087F0000003E4140413E000040407E41417E0000",
            INIT_RAM_39 => X"00013F4141410000033E4141414100000041413E41410000083E4949493E0000",
            INIT_RAM_3A => X"0079457941410000007E417E40C00000033E494949490000003F494949490000",
            INIT_RAM_3B => X"00413F41413F0000004E5171514E0000003E410F413E0000007E417E40400000",
            INIT_RAM_3C => X"0C18306030180C0030180C060C183000007C0010107C101000FE00FE00FE0000",
            INIT_RAM_3D => X"0000DC7600DC76001818007E0018180070D8D8181818181818181818181B1B0E",
            INIT_RAM_3E => X"103868CC0406020300000018000000000000001818000000000000386C6C3800",
            INIT_RAM_3F => X"007E42000000000000007C7C7C7C000000000078201048303C4299A1A199423C"
        )
        port map (
            DO => prom_inst_0_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => prom_inst_0_AD_i
        );

end Behavioral; --Gowin_pROM_font
